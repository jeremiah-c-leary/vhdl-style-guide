
architecture RTL of FIFO is

begin

  process
  begin

    LOOP_LABEL : loop

    end loop;

    -- Violations below

    LOOP_LABEL : loop

    end loop;

  end process;

end;
