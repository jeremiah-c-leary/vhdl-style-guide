
entity FIFO is

end entity;

entity FIFO is

end entity;

entity FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MYFIFO is

end entity;

entity MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity MYFIFP is

end entity;

entity MYFIFO is

end entity;

entity E_MYFIFO_A is

end entity;

entity E_MYFIFO_A is

end entity;

entity MYFIFO_A is

end entity;

entity MYFIFO_A is

end entity;

