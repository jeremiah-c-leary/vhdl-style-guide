
entity FIFO is

end entity FIFO;


entity FIFO is

end entity FIFO;


entity FIFO2 is

end entity FIFO2;
