
architecture rtl of fifo is

  constant width  : integer := 32;
  signal   height : integer := 4;

  constant width  : integer := 32;
  constant height : integer := 4;

begin

end architecture rtl;
