
library IEEE;

library IEEE;
