
architecture rtl of fifo is

begin

  GEN_LABEL : for x in range (3 downto 0) GENERATE

  end generate;

  GEN_LABEL : for x in range (3 downto 0) GENERATE

  end GENERATE;

end architecture;
