
architecture RTL of FIFO is

begin

  block_label_blk : block is begin end block block_label_blk;

  block_label : block is begin end block block_label;

end architecture RTL;
