
entity entity1 is
  port (
    port1 : in    std_logic;
    port2 : out   std_logic;
    port3 : inout std_logic;
    port4 : in    std_logic;
    port5 : out   std_logic;
    port6 : inout std_logic
  );
end entity entity1;

architecture arch of entity1 is

begin

end architecture arch;
