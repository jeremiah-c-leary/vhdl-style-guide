
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--+-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--!-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--+--------------------------------[ abcdef ]===================================
-- Comment
--------------------------------------------------------------------------------

--+-[ abcdef ]==================================================================
-- Comment
--------------------------------------------------------------------------------

--+------------------------------------------------------------------[ abcdef ]=
-- Comment
--------------------------------------------------------------------------------
architecture rtl of fifo is

  --+-------------------------------[ abcdef ]==================================
  -- Comment
  ------------------------------------------------------------------------------

  signal sig1 : std_logic;

begin

end architecture rtl;
-- comment
-- comment

--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

architecture rtl of FIFO is

begin

    inst_dummy : entity lib.module
    port map (
      -- Clocks
      clk   => clk
      --
      -- Dummy comment
      --
      data_i => data_i
    );

end architecture rtl;
