
architecture RTL of FIFO is

  procedure PROC1 is begin end procedure proc1;

  PROCEDURE PROC1 IS BEGIN END PROCEDURE PROC1;

begin

end architecture RTL;
