
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  COMPONENT fifo is--Some Comemnt
   -- Some COmment

  end component fifo;

  Component fifo is--Other comment
  -- Some Comment
 

  end component fifo;

begin

end architecture RTL;
