
architecture rtl of fifo is

begin

  process begin

    report "hello" severity FAILURE;

    report "hello"
      severity FAILURE;

  end process;

end architecture rtl;
