
architecture RTl of FIFO is

  component fifo

  end component fifo;

  -- Failures below

  component fifo

  end component fifo;

begin

end architecture RTL;
