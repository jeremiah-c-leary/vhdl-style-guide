
architecture rtl of fifo is

begin

  process
  begin
    case expression is
      when OTHERS =>

    end case;

    case expression is
      when OTHERS =>

    end case;
  end process;

end architecture;
