
architecture RTL of FIFO is

  procedure proc_name (
    constant a : in integer;
    signal b : in std_logic;
    variable c : in std_logic_vector(3 downto 0);
    signal d : out std_logic) is
    constant con1 : integer := 0;
    variable var1 : integer := 12;
    use ieee.std_logic_1164.all;
  begin
  end procedure proc_name;

  procedure proc_name (
      constant a : in integer;
     signal b : in std_logic;
    variable c : in std_logic_vector(3 downto 0);
signal d : out std_logic) is
    constant con1 : integer := 0;
    variable var1 : integer := 12;
    use ieee.std_logic_1164.all;
    
  begin
  end procedure proc_name;

  procedure proc_name (
constant a : in integer;
      signal b : in std_logic;
     variable c : in std_logic_vector(3 downto 0);
    signal d : out std_logic) is
    constant con1 : integer := 0;
    variable var1 : integer := 12;
    use ieee.std_logic_1164.all;
    
  begin
  end procedure proc_name;

begin

end architecture RTL;
