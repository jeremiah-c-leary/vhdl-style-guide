
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo is

end component fifo;

  component fifo is

    end component fifo;

begin

end architecture RTL;
