
architecture RTL of FIFO is

  signal sig1 : std_logic_vector(3 downto 0);

  signal sig1 : std_logic_vector(3 downto 0   );

begin

  a <= (b or ((c and d and e)));
  a <= (b or ((c and d and e))
       );
  a <= (b or ((c and d and e))
);

  a <= (b or ((c and d and e  )  )  );

  a <= (b or ' ');
  a <= (b or ' ' );

end architecture RTL;
