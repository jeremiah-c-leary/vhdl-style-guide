
architecture RTL of FIFO is

begin


  process 
  begin
  END process;

  -- Violations below

  process 
  begin
  END process;

end architecture RTL;
