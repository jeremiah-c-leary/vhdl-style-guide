
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo is

  end component FIFO;

  component fifo is

  end component Fifo;

begin

end architecture RTL;
