
architecture rtl of fifo is

  signal   width  : integer := 32;

  constant height : integer := 4;

  signal   width  : integer := 32;
  signal   height : integer := 4;

begin

end architecture rtl;
