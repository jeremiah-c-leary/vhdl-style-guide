
entity FIFO is end entity;
entity E_FIFO is end entity;
entity FIFO_A is end entity;
entity E_FIFO_A is end entity;

entity FIFO is end entity;
entity E_FIFO is end entity;
entity FIFO_A is end entity;
entity E_FIFO_A is end entity;

entity FIFO is end entity;
entity E_FIFO is end entity;
entity FIFO_A is end entity;
entity E_FIFO_A is end entity;

entity FIFO is end entity;
entity E_FIFO is end entity;
entity FIFO_A is end entity;
entity E_FIFO_A is end entity;

entity MY_FIFO is end entity;
entity E_MY_FIFO is end entity;
entity MY_FIFO_A is end entity;
entity E_MY_FIFO_A is end entity;

entity MY_FIFO is end entity;
entity E_MY_FIFO is end entity;
entity MY_FIFO_A is end entity;
entity E_MY_FIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

entity MYFIFO is end entity;
entity E_MYFIFO is end entity;
entity MYFIFO_A is end entity;
entity E_MYFIFO_A is end entity;

-- Test Pascal_Snake_Case

entity MYFIFO_GREENRED_BLUE is end entity;
entity E_MYFIFO_GREENRED_BLUE is end entity;
entity MYFIFO_GREENRED_BLUE_A is end entity;
entity E_MYFIFO_GREENRED_BLUE_A is end entity;

entity MY_FIFO_GREEN_RED_BLUE is end entity;
entity E_MY_FIFO_GREEN_RED_BLUE is end entity;
entity MY_FIFO_GREEN_RED_BLUE_A is end entity;
entity E_MY_FIFO_GREEN_RED_BLUE_A is end entity;

-- Test RelaxedPascalCase

entity MYFIFO is end entity;
entity MYFIFO is end entity;
entity MYFIFO is end entity;
entity MYFIFO is end entity;
entity MYFIFO is end entity;
entity MYFIFO is end entity;
entity MYFIFO is end entity;
