

architecture ARCH of ENTITY is

  signal a_sig : std_logic_vector(31 downto 0);
   signal a_SIg :  std_logic_vector(31 downto 0);
  Signal b_sig: std_logic_vector(31 downto 0);
 signal  b_sig : std_logic_vector(31 downto 0);
  signal  siG : std_logic_vector(31 downto 0);
  signal d_sig :std_logic_vector(31 downto 0);
  siGNal e_sig: std_logic_vector(31 downto 0) := "0";
  signal   SIg : STD_LOGIC_VECTOR(31 downto 0);
  signAL sig :   std_logic_vector(GENERIC_1 downto 0);
  signal sig :std_logic_vector(31 downto 0);
     signal sIg : std_logic_vector(31 downto 0);
  signal sig :   STD_LOGIC_VECTOR (31 downto 0) := (others => '0');

  signal e_sig1, d_sig2 : std_logic;
  signal a_sig10, c_sig2: std_logic;
  signal b_sig100, b_sig2 :std_logic_vector (31 downto 0);
  signal c_sig1000, a_sig2:std_logic;
  
  signal w_sig1 : t_User_Defined_Type;

begin

end architecture ARCH;
