
architecture RTL of FIFO is

  shared variable c_width : integer := 16;
  shared    variable c_depth : integer := 512;

begin

end architecture RTL;
