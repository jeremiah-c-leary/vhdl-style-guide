
architecture rtl of fifo is

  file defaultimage : load_file_type open READ_MODE is load_file_name;
  file defaultimage : load_file_type open WRITE_MODE is load_file_name;
  file defaultimage : load_file_type open APPEND_MODE is load_file_name;

  file defaultimage : load_file_type open READ_MODE is load_file_name;
  file defaultimage : load_file_type open WRITE_MODE is load_file_name;
  file defaultimage : load_file_type open APPEND_MODE is load_file_name;

  file defaultimage : load_file_type open READ_MODE is load_file_name;
  file defaultimage : load_file_type open WRITE_MODE is load_file_name;
  file defaultimage : load_file_type open APPEND_MODE is load_file_name;

begin

end;
