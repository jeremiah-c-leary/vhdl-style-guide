
architecture rtl of fifo is

begin

  x <= a and b or c nand d nor e xor f xnor g;

  x <= a and b or c nand d nor e xor f xnor g;

end architecture;
