
architecture RTL of FIFO is

begin

  process
  begin

    label : for index in 4 to 23 loop

    end loop;

    loop_label : for index in 4 to 23 loop

    end loop;

  end process;

end;
