
--This should pass
context c1 is

end context c1;

--These should fail
CONTEXT c1 is
end context c1;

CoNtExT c1 is

end context c1;
