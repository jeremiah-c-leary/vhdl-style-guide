
package fifo_pkg is

  signal wr_en        : std_logic;
  signal rd_en        : std_logic;
  constant c_constant : integer;

  signal wr_en : std_logic;
  signal rd_en   : std_logic;
  constant c_constant : integer;

end package;

