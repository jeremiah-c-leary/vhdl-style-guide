
architecture RTL of FIFO is

begin

  process 
  begin
  end process;

  process 
  begin
  end postponed process;

  -- Violations below

  process 
  begin
  end    process;

  process 
  begin
  end    postponed process;

end architecture RTL;
