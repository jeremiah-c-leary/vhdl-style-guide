
architecture rtl of fifo is

begin

  process begin

    REPORT "hello";

    report "hello";

  end process;

end architecture rtl;
