
--------------------------------------------------------------------------------
-- Comment
-- Comment
-- Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--+ Comment
--+ Comment
--+ Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--| Comment
--| Comment
--| Comment
--| Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--!-- Comment
--!-- Comment
--!-- Comment
--!-- Comment
--------------------------------------------------------------------------------

-- comment
-- comment
-- comment
-- comment
-- comment


--+ Comment
--+ Comment
--+ Comment


--| Comment
--| Comment
--| Comment
--| Comment

  ------------------------------------------------------------------------------
  --+ Comment
  --+ Comment
  --+ Comment
  ------------------------------------------------------------------------------

architecture rtl of FIFO is

begin

    inst_dummy : entity lib.module
    port map (
      -- Clocks
      clk   => clk
      --
      -- Dummy comment
      --
      data_i => data_i
    );


    -- Comment

end architecture rtl;

