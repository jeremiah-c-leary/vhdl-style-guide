
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--+-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--!-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--!---------------------------------[ abcdef ]==================================

--------------------------------------------------------------------------------
-- Comment
--!-[ abcdef ]==================================================================

--------------------------------------------------------------------------------
-- Comment
--!------------------------------------------------------------------[ abcdef ]=

-- comment
-- comment
