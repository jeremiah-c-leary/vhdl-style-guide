
architecture RTl of FIFO is

  component fifo is

  end COMPONENT fifo;

  -- Failures below

  component fifo is

  end COMPONENT fifo;

  component fifo is

  end COMPONENT fifo;

begin

end architecture RTL;
