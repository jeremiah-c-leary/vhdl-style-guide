

package PACK1 is

end package PACK1;

package PACK2 is

end package;

package PACK3 is

end;

