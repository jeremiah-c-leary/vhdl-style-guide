
architecture rtl of fifo is

begin

  x <= a and b or c nand d nor e xor f xnor g;

  x <= a AND b OR c NAND d NOR e XOR f XNOR g;

end architecture;
