
architecture RTL of FIFO is

  constant c_width : integer := 16;
  constant c_depth : integer := 512;
  constant c_word : integer := (12, 13, 15);

begin

  process

    constant c_width : integer :=    16;
    constant c_depth : integer :=512;
    constant c_word : integer :=(12, 13, 15);
    constant c_word : integer :=          (12, 13, 15);

  begin end process;

end architecture RTL;
