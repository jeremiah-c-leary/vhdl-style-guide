
library ieee;

library IEEE;

