
architecture RTL of FIFO is

begin

  process
  begin

    for_label : for index in 4 to 23 loop

    end loop for_label;

    FOR_LABEL : for index in 4 to 23 loop

    end loop FOR_LABEL;

    For_label : for index in 4 to 23 loop

    end loop For_label;

  end process;

end;
