
architecture rtl of fifo is

  alias designator is name;

  alias designator is name;

begin

end architecture rtl;
