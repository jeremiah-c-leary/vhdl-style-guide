

architecture ARCH of ENTITY is

  variable a_sig : std_logic_vector(31 downto 0);
   variable a_SIg :  std_logic_vector(31 downto 0);
  Variable b_sig: std_logic_vector(31 downto 0);
 variable  b_sig : std_logic_vector(31 downto 0);
  variable  siG : std_logic_vector(31 downto 0);
  variable d_sig :std_logic_vector(31 downto 0);
  varIAble e_sig: std_logic_vector(31 downto 0) := "0";
  variable   SIg : STD_LOGIC_VECTOR(31 downto 0);
  variabLE sig :   std_logic_vector(GENERIC_1 downto 0);
  variable sig :std_logic_vector(31 downto 0);
     variable sIg : std_logic_vector(31 downto 0);
  variable sig :   std_logic_vector(31 downto 0) := (others => '0');

  variable e_sig1, d_sig2 : std_logic;
  variable a_sig1, c_sig2: std_logic;
  variable b_sig1, b_sig2 :std_logic;
  variable c_sig1, a_sig2:std_logic;

begin

end architecture ARCH;
