
architecture rtl of ENT is
begin
end RTL;

architecture rtl of ENT is
begin
end rtl;

architecture rtl of ENT is
begin
end Rtl;

architecture rtl of ENT is
begin
end;

architecture rtl of ENT is
begin
end architecture;
