
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    target := expression;

    target(i) := expression;

    ( element_association ) := expression;

    ( element_association, element_association, element_association ) := expression;

  end process;

end architecture RTL;
