architecture RTL of FIFO is
constant fifo_wr : std_logic;

constant fifo_wr : std_logic_vector(3 downto 0);

constant fifo_wr : std_logic_vector(3 downto 0) := "000";

constant fifo_wr, fifo_rd, fifo_empty : std_logic := '1';

constant
fifo_wr
,
fifo_rd
,
fifo_empty
:
std_logic
:=
'1'
;

constant
fifo_wr
,
fifo_rd
,
fifo_empty
:
std_logic_vector( 3 downto 0 )
:=
'1'
;

begin

end architecture RTL;
