
entity FIFO is

end entity FIFO;

entity FIFO is

end entity;

entity FIFO is

end;

entity FIFO is

end FIFO;
