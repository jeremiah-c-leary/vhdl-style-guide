
architecture rtl of fifo is

begin

  process begin

    loop end loop;

    LOOP END LOOP;

  end process;

end;
