
package fifo_pkg is

end package;

package fifo_pkg is --comment


end package;
