
library ieee;
	--Comment
  use ieee.std_logic_1164.all;
	--Comment
  use ieee.numeric_std.all;

library ieee;
	-- Comment
  use ieee.std_logic_1164.all;
	-- Comment
	-- Comment 2
	-- Comment 3
  use ieee.numeric_std.all;
	-- Comment
  use ieee.std_logic_arith.all;

library ieee;
	-- Comment
	use ieee.std_logic_1164.all;

