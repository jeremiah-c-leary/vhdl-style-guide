
architecture RTL of ENT is begin end architecture RTL;

architecture RTL of ENT is

begin
end;

architecture RTL of ENT is
-- Some domment

begin
end;

architecture RTL of ENT is--some comment

begin
end;

