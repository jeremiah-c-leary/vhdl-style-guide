
architecture RTl of FIFO is

  component FIFO is

  end component fifo;

  -- Failures below

  component FIFO is

  end component fifo;

  component FIFO is

  end component fifo;

begin

end architecture RTL;
