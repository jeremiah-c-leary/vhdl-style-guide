
architecture rtl of fifo is

begin

  process begin

    while (condition) loop end loop;

    while (condition) loop end loop;

    while condition loop end loop;

  end process;

end;
