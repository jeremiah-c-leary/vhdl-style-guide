
architecture rtl of fifo is

  procedure proc is
  begin
  end procedure proc;

  procedure proc is
  begin
  end procedure proc;

  function func return integer is
  begin
  end function func;

  function func return integer is
  begin
  end func;

  procedure proc;

  function func return integer is
  begin
  end func;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end procedure proc;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end procedure proc;

begin

end architecture rtl;
