
architecture rtl of fifo is

  type t_record is record
  end record;

  type t_record is
  record end record;

begin

end architecture rtl;
