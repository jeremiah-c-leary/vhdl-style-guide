
architecture ARCH of ENTITY_1 is

  function func_1 (a : integer; b : integer;
             c : unsigned(3 downto 0);
     d : std_logic_vector(7 downto 0);
        e : std_logic) return integer is
  begin

  end;

begin


end architecture ARCH;
