
architecture rtl of fifo is

begin

  x <= a SLL b SRL c SLA d SRA e ROL f ROR g;

  x <= a SLL b SRL c SLA d SRA e ROL f ROR g;

end architecture;
