
package my_pkg is NEW my_generic_pkg
  generic map (
    g_my_generic => 2
  );

package my_pkg is NEW my_generic_pkg
  generic map (
    g_my_generic => 2
  );
