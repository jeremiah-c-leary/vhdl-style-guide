
entity fifo is

end entity;

entity FIFO is

end entity;

entity Fifo is

end entity;

entity MY_FIFO is

end entity;

entity my_fifo is

end entity;

entity MyFifo is

end entity;

entity myFifo is

end entity;

