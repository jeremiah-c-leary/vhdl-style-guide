
architecture rtl of fifo is

  type integer_file is file OF integer;

  type integer_file is file OF integer;

  type integer_file is file OF integer;

begin

end;
