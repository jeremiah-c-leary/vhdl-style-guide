
architecture rtl of fifo is

  component my_block is
  end component;

  -- synthesis translate_off

  component my_block is
  end component;

  -- synthesis translate_off

begin

end architecture;
