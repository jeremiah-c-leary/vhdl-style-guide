
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component FIFO is

  end component fifo;

  component Fifo is

  end component fifo;

begin

end architecture RTL;
