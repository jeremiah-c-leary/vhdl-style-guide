
architecture RTL of ENTITY1 is

  procedure AVERAGE_SAMPLES (
    constant a : in integer;
    signal d : out std_logic
  );

begin

  PROC1 : process () is
  begin

    Average_samples();

  end process PROC1;

end architecture RTL; 

