
entity FIFO is

end entity fifo;

entity FIFO is

end entity FIFO;

entity FIFO is

end entity Fifo;

