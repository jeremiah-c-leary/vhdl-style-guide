-- ANSI "���" comment
