
entity FIFO is

end entity;


entity FIFO is --Comment
--Comment
--Comment


end entity;
