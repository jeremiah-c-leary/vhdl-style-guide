
architecture rtl of fifo is

begin

  process begin

    REPORT "hello";

    REPORT "hello";

  end process;

end architecture rtl;
