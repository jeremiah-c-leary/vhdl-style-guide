
entity FIFO is

end ENTITY fifo;

entity FIFO is

end ENTITY FIFO;

entity FIFO is

end ENTITY FIFO;

