
architecture RTL of FIFO is

  function func1 return integer is begin END function func1;

  function func1 return integer is begin END function func1;

  function func1 return integer is begin END function func1;

begin

end architecture RTL;
