
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo is

  end component fifo;

  signal sig1 : std_logic;

begin

end architecture RTL;
