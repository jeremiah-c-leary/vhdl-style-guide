
entity FIFO is

end entity FIFO;

--vhdl_comp_off
entity FIFO is
--vhdl_comp_on

entity FIFO is

end entity;
