
architecture rtl of fifo is

  type t_record is
  record
    a : std_logic;
    b : std_logic;
  end record t_record;

  type t_record is
  record
    a : std_logic;
    b : std_logic;
  end record t_record;

  type t_record is
  record
    a : std_logic;
    b : std_logic;
  end record t_record;

  type t_record is record a : std_logic; b : std_logic; end record;

  type t_record is record
    a : std_logic;
    b : std_logic;
  end record t_record;

begin

end architecture rtl;
