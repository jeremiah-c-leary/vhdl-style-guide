
architecture RTL of FIFO is

  constant c_width : integer := 16;

  constant c_depth : integer
  := 512;

begin

end architecture RTL;
