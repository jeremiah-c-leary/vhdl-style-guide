

library lib1
-- Comment 1
  use lib1.all

library lib1
  -- Comment 1
  use lib1.all

