entity FIFO is
generic ( );
end entity FIFO;

entity FIFO is
generic (

);
end entity FIFO;

entity FIFO is
generic
(
)
;
end entity FIFO;
