
architecture RTL of FIFO is

begin


  process is
  begin
  end process;

  process (a, b) is
  begin
  end process;

  -- Violations below

  process is
  begin
  end process;

  process (a, b)is
  begin
  end process;

  process(a,b)is begin end process;

end architecture RTL;
