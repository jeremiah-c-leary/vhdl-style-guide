

architecture ARCH of ENTITY1 is

  signal sig1 : std_logic;
  file fil1 : something...;
  -- Comment1
  type typ1 : fifo_sigs;
  subtype sub1 : other_type;
  -- Comment1
  variable var1 : integer;
  constant con1 : integer := 0;

  attribute att1 : some_attr;

begin

end architecture ARCH;
