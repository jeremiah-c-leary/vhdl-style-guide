
architecture RTL of FIFO is

  attribute max_delay : time;

  ATTRIBUTE MAX_DELAY : TIME;

begin

end architecture RTL;
