
package body test is

  type flag_pt is protected body
  END protected body;

  type flag_pt is protected body
  END protected body;

end package body test;

architecture rtl of test is

  type flag_pt is protected body
  END protected body;

  type flag_pt is protected body
  END protected body;

begin

end architecture rtl;
