
context c1;

context c2;

context c2;
