
entity FIFO is

end entity;


entity --Comment
--Comment
--Comment
FIFO is

end entity;
