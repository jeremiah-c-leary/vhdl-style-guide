
architecture rtl of fifo is

begin

  process begin

    loop end loop;

    LOOP END loop;

  end process;

end;
