
entity FIFO is
  port (
    I_INPUT : in integer;
    O_OUTPUT : out integer
  );
end entity FIFO;

entity FIFO is
  port (
    I_INPUT : in integer;
    O_OUTPUT : out integer
  );
end entity FIFO;

entity FIFO is
  generic (
    G_GENERIC : integer
  );
  port (
    I_INPUT : in integer;
    O_OUTPUT : out integer
  );
end entity FIFO;
