
architecture RTL of FIFO is

begin


  process
  BEGIN
  end process;

  -- Violations below

  process
  BEGIN
  end process;

end architecture RTL;
