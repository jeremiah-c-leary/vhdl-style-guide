
architecture rtl of fifo is

begin

  x <= a sll b srl c sla d sra e rol f ror g;

  x <= a SLL b SRL c SLA d SRA e ROL f ROR g;

end architecture;
