

use ieee.std_logic_1164.all;

use my_lib, otherlib.my_math_stuff.multiply;

use yetanotherlib.std_logic;

