
architecture RTL of ENTITY1 is

  subtype st_range is range 0 to 9;
  subtype st_width is range 16 to 128;

  subtype subt_range is range 0 to 9;
  subtype subt_width is range 16 to 128;

  subtype stRange is range 0 to 9;
  subtype stWidth is range 16 to 128;

begin

end architecture RTL;

