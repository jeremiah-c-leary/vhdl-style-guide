
entity FIFO is
  port (
    I_INPUT : in std_logic
  );
begin
end entity;


entity FIFO is
  port (
    I_INPUT : in std_logic
  );
begin
end entity;

