
entity FIFO is
  port (
    port1 : in std_logic
  );
end entity;

entity FIFO is
  port (
    port1 : in std_logic
  );

end entity;

entity FIFO is
  port (
    port1 : in std_logic
  );





end entity;
