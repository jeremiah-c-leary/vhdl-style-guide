
architecture RTL of FIFO is

  procedure proc_name (
    constant a : in integer;
    signal b : in std_logic;
    variable c : in std_logic_vector(3 downto 0);
    signal d : out std_logic) is
  begin
  end procedure proc_name;

begin

  proc_Name (0, '1', x"00", sig1);

  PROC_NAME (0, '1', x"00", sig1);

end architecture RTL;
