
entity FIFO is
begin
end entity;

entity FIFO is
BEGIN
end entity;

