

architecture ARCH of ENT is

  signal sig1 : std_logic;
  signal sig2 : std_logic;;
  signal sig3 : std_logic;;;

  signal sig4 : std_logic;signal sig5 : std_logic;;;

  signal sig6 : std_logic;;signal sig7 : std_logic;signal sig8 : std_logic;;;

  signal sig9 : std_logic;;;signal sig10 : std_logic;;signal sig11 : std_logic;;;

  signal sig12 : std_logic;signal sig13 : std_logic;signal sig14 : std_logic;

  -- Checking comments are ignored
  signal sig15 : std_logic;signal sig16 : std_logic;signal sig17 : std_logic; --;;;


  signal sig18 : std_logic;;;signal sig19 : std_logic;;signal sig20 : std_logic;;; --;;;

begin

end architecture ARCH;
