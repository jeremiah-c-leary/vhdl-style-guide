
architecture rtl of fifo is

  constant cons1 : t_type :=
 (
    1 => func1(std_logic_vector(G_GEN), G_GEN2),
 2 => func1(std_logic_vector(G_GEN3), G_GEN4)
 );

begin

end architecture rtl;
