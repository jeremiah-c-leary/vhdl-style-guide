
--This should pass
context c1 is

end context c1;

context c1 is
end context c1;

context c1 is
-- Comment
end context c1;
