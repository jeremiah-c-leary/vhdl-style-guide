
entity fifo is

end entity;

entity FIFO is

end entity;

entity Fifo is

end entity;

entity MY_FIFO is

end entity;

entity my_fifo is

end entity;

entity MyFifo is

end entity;

entity myFifo is

end entity;

entity e_myFifo is

end entity;

entity e_MyFifo is

end entity;

entity e_MyFIFo is

end entity;

entity e_myFIFo is

end entity;

entity MyFIFp is

end entity;

entity myFIFo is

end entity;

entity e_MyFIFo_a is

end entity;

entity e_myFIFo_a is

end entity;

entity MyFIFo_a is

end entity;

entity myFIFo_a is

end entity;

