
architecture RTl of FIFO is

  COMPONENT fifo is

  end component fifo;

  -- Failures below

  COMPONENT fifo is

  end component fifo;

  COMPONENT fifo is

  end component fifo;

begin

end architecture RTL;
