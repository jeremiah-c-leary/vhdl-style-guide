
architecture RTL of FIFO is begin end architecture RTL;

architecture RTL of FIFO is
begin
end architecture RTL;

-- This should fail

  architecture RTL of FIFO is

     begin

end architecture RTL;
