
library ieee;

LIBRARY ieee;
