
architecture RTL of FIFO is

begin


  PROC_LABEL : process
  begin
  end process;

  process
  begin
  end process;

  -- Violations below

  
  PROC_LABEL : process (b) is
  begin
  end process;

  




  PROC_LABEL : process (c) is
  begin
  end process;

end architecture RTL;
