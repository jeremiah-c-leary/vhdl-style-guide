

architecture Arch of ENTITY is

begin

End  architecture ARCH;

  architecture ARCH of EntITY is

begin

end Architecture;
architecture  ARCH  of  ENTITY  is

begin

end  architecture ARCH

 Architecture ARch Of entity Is

 begin

 eND architecture ArCh

architecture ARch
 of ENTITY is

BEGIN

 end archITecture   ARCH

architecture ARCH of ENTITY iS
begin
end architecture ARCH;

architecture ARCH of ENTITY is

begin

  process () is
  begin
  end process;

end architecture ARCH;

architecture ARCH of ENTITY is

begin

  process () is
  begin
  end process;

end ARCH;

-- Comment

architecture ARCH of ENTITY is

begin

  GEN1 : if CONDITION = 1 generate

    process () is
    begin
    end process;

  end generate;

  END_PROC : process () is
    begin
    end process END_PROC;

  end_signal <= '0';

end;

-- Comment

architecture ARCH of arch is

begin

end architecture ARCH;
