
package pkg is

  procedure my_proc is new MY_GENERIC_PROC
    generic map (
      test => 2
    );

  function my_func is new MY_GENERIC_FUNC
    generic map (
      test => 2
    );

  procedure my_proc is new MY_GENERIC_PROC
    generic map (
      test => 2
    );

  function my_func is new MY_GENERIC_FUNC
    generic map (
      test => 2
    );

  procedure my_proc is new MY_GENERIC_PROC
    generic map (
      test => 2
    );

  function my_func is new MY_GENERIC_FUNC
    generic map (
      test => 2
    );

end package;
