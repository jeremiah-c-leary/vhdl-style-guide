
entity FIFO is

end entity fifo;

entity FIFO is

end entity fifo;

entity FIFO is

end entity fifo;

