
package fifo_pkg is

end package;

package fifo is

end package;

