package test is

  type flag_pt is protected
  end protected;

  type flag_pt is protected
  END protected;

end package test;

architecture rtl of test is

  type flag_pt is protected
  end protected;

  type flag_pt is protected
  END protected;

begin

end architecture rtl;
