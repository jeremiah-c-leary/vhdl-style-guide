
package fifo_pkg is

end package;

PACKAGE fifo_pkg is

end package;

