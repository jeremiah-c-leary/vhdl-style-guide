
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block is
  begin
    a <= b;

  end block;

  BLOCK_LABEL : block is
  begin
    a <= b;
  end block;

end architecture RTL;
