
architecture RTl of FIFO is

  component fifo IS

  end component fifo;

  -- Failures below

  component fifo IS

  end component fifo;

  component fifo IS

  end component fifo;

begin

end architecture RTL;
