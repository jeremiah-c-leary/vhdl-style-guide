
architecture RTL of FIFO is

  subtype state_machine is subtype_indication;

  -- Violations below

  subtype state_machine is subtype_indication;

begin

end architecture RTL;
