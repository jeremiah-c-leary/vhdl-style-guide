
architecture rtl of fifo is

begin

  block_label : block is
  begin

  end block block_label;

      ------------------------------<-    80 chars    ->------------------------------
  --! FPGA RX to Avalon-ST TX interface
 --------------------------------------------------------------------------------

  ------------------------------<-    80 chars    ->------------------------------
  --------------------------------------------------------------------------------

  ------------------------------<-    80 chars    ->------------------------------

    ------------------------------<-    80 chars    ->------------------------------
      --! FPGA RX to Avalon-ST TX interface
  --! FPGA RX to Avalon-ST TX interface
     --! FPGA RX to Avalon-ST TX interface
  --------------------------------------------------------------------------------

  ------------------------------<-    80 chars    ->------------------------------
    --! FPGA RX to Avalon-ST TX interface
  --! FPGA RX to Avalon-ST TX interface
    --! FPGA RX to Avalon-ST TX interface
   --! FPGA RX to Avalon-ST TX interface
       --------------------------------------------------------------------------------

  -- vsg_off comment_010
  ------------------------------<-    80 chars    ->------------------------------
    --! FPGA RX to Avalon-ST TX interface
  --! FPGA RX to Avalon-ST TX interface
    --! FPGA RX to Avalon-ST TX interface
   --! FPGA RX to Avalon-ST TX interface
       --------------------------------------------------------------------------------
  -- vsg_on comment_010

  -- vsg_off signal_001
         ------------------------------<-    80 chars    ->------------------------------
     --! FPGA RX to Avalon-ST TX interface
 --------------------------------------------------------------------------------
  -- vsg_on signal_001

  -- vsg_off signal_001
------------------------------<-    80 chars    ->------------------------------
      --------------------------------------------------------------------------------
  -- vsg_on signal_001

  a <= b;

end architecture rtl;
