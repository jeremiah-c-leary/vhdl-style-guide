-------------------------------------------------------------------------------
--  Next line is a failure
-------------------------------------------------------------------------------

architecture RTL of ENT is

  signal a : std_logic;

  signal a : std_logic_vector(15 downto 0);

begin

end architecture RTL;
