
package fifo_pkg is

END package;

package fifo_pkg is

END package;
