
#ifdef G_I2C_ENABLE

 #ifdef G_I2C ENABLE
