entity FIFO is
port ( );
end entity FIFO;

entity FIFO is
port (

);
end entity FIFO;

entity FIFO is
port
(
)
;
end entity FIFO;
