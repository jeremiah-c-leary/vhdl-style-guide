
entity entity1 is
  port (
    i_port1 : in    std_logic;
    i_port2 : in    std_logic;

    o_port3 : out   std_logic;
    o_port4 : out   std_logic
  );
end entity;
