
configuration CFG of FIFO is
end configuration CFG;


configuration CFG of FIFO is
end;


configuration CFG of FIFO is
end configuration;


configuration CFG of FIFO is
end CFG;

