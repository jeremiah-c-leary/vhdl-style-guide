
entity FIFO is

end entity FIFO;

--vhdl_comp_off
entity FIFO is
--vhdl_comp_on

entity FIFO is

-- synthesis
-- synthesis something
-- synthesis something else
-- synthesis something else entirely

-- pragma
-- pragma something
-- pragma something else
-- pragma something else entirely

-- altera
-- altera something
-- altera something else
-- altera something else entirely

-- RTL_SYNTHESIS
-- RTL_SYNTHESIS ON
-- RTL_SYNTHESIS OFF
-- RTL_SYNTHESIS something

-- synopsys 
-- synopsys something
-- synopsys something else
-- synopsys something else entirely

-- xilinx 
-- xilinx something
-- xilinx something else
-- xilinx something else entirely

end entity;
