
architecture RTL of FIFO is

begin


  PROC_LABEL : process is
  begin
  end process;

  -- Violations below

  proc_label : process is
  begin
  end process;

end architecture RTL;
