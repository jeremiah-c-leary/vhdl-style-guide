
architecture RTL of ENT is
begin
end RTL;

architecture rtl of ENT is
begin
end rtl;

architecture Rtl of ENT is
begin
end Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;
