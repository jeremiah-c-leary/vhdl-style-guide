
architecture ARCH of ENTITY is

  signal sig1 : std_logic;        -- comment
  signal sig1 : std_logic;    -- comment
  signal sig1 : std_logic;  -- comment
  signal sig1 : std_logic;         -- comment
  signal sig1 : std_logic; -- comment

begin

end architecture ARCH;
