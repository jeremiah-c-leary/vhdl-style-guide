
package body fifo_pkg is

end package body fifo_pkg;

package body fifo_pkg is

end package body fifo_pkg;

package body fifo_pkg is

end package body;

