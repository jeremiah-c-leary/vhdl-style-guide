
architecture rtl of fifo is

  file defaultimage : load_file_type open read_mode is load_file_name;
  file defaultimage : load_file_type open write_mode is load_file_name;
  file defaultimage : load_file_type open append_mode is load_file_name;

  file defaultimage : load_file_type open READ_MODE is load_file_name;
  file defaultimage : load_file_type open WRITE_MODE is load_file_name;
  file defaultimage : load_file_type open APPEND_MODE is load_file_name;

  file defaultimage : load_file_type open Read_Mode is load_file_name;
  file defaultimage : load_file_type open Write_Mode is load_file_name;
  file defaultimage : load_file_type open Append_Mode is load_file_name;

begin

end;
