

architecture RTL of ENT is

begin

  -- vsg-disable-next-line process_016
  process (A) is
  begin
    -- vsg-disable-next-line process_018
  end process;

  process (A) is
  begin
  end process;

  -- vsg-disable-next-line process_016
  -- vsg-disable-next-line process_002
  process(A)is
  begin

  -- vsg-disable-next-line process_018
  end process;

  process (A) is
  begin
  end process;

  -- vsg-disable-next-line architecture_024
end architecture;
