
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    PROC_LABEL : proc(a, b, c);

    PROC_LABEL : proc;

    proc(a, b, c);

    proc(x"1", d"5", o"X");

    proc;

  end process;

end architecture RTL;
