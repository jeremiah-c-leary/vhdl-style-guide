
architecture rtl of fifo is

begin

  PROC_LABEL : postponed process begin end process;

  PROC_LABEL : postponed -- Comment
  process begin end process;

  PROC_LABEL : postponed -- Comment




  process begin end process;

end;
