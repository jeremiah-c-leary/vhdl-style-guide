
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  component fifo is

  end component;

begin

end architecture RTL;
