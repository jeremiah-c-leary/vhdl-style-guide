
architecture rtl of fifo is

  alias designator is name;

  signal sig1 : std_logic;alias designator is name;

  signal sig1 : std_logic; alias designator is name;

begin

end architecture rtl;
