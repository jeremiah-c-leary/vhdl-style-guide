
architecture RTL of FIFO is

  subtype state_machine IS subtype_indication;

  -- Violations below

  subtype state_machine IS subtype_indication;

begin

end architecture RTL;
