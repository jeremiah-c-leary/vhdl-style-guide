
architecture rtl of fifo is

begin

  process begin

    for x in (31 downto 0) loop end loop;

    for X in (31 downto 0) loop end loop;

  end process;

end;
