
architecture RTL of FIFO is

  procedure proc1 is
  begin

  end procedure proc1;

  -- Fixes follow

  procedure proc1 is
  begin
  end procedure proc1;

begin

end architecture RTL;
