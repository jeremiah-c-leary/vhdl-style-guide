
architecture RTL of ENTITY1 is


begin

  PROC_NAME : process () is

    variable var1 : std_logic;
    variable var2 : std_logic;
    variable var3 : std_logic;
    variable var4 : std_logic;

  begin

    Var1 <= '0';

    if (VAR2 = '0') then
      vaR3 <= '1';
    elsif (var2 = '1') then
      VAR4 <= '0';
    end if;

    vaR1 <= VAR2 & Var3 & vAr4;

  end process PROC_NAME;

end architecture RTL;

