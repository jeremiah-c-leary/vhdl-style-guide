library ieee;

package body fifo_pkg is

end package body;

-- Violation below

package body fifo_pkg is

end package body;
-- Comments could be allowed


library ieee;
package body fifo_pkg is

end package body;
entity fifo is

end entity fifo;
