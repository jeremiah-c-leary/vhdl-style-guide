
architecture RTL of FIFO is

  attribute  coordinate  of  comp_1:component is  (0.0, 17.5);

  -- Violations below

  attribute  coordinate  of  comp_1:component is  (0.0, 17.5);

begin

end architecture RTL;
