
entity ENTITY1 is
  port (PORT_1 : in std_logic_vector(12 downto 0),
    PORT_2 : out std_logic_vector(0 to 25)
  );
end entity ENTITY1;

