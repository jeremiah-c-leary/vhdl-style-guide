
architecture RTL of ENT is
begin
end architecture RTL;

architecture RTL of ENT is
begin
end architecture RTL;

architecture RTL of ENT is
begin
end architecture;

architecture RTL of ENT is
begin
end architecture;

architecture RTL of ENT is
begin
end architecture
;

architecture RTL of ENT is
begin
end architecture--Comment
;
