
LABEL : assert TRUE
  report "This is a string"
  severity WARNING;


assert TRUE
  report "This is a string"
  severity WARNING;

LABEL : assert TRUE
  report "This is a string";

LABEL : assert TRUE
  severity WARNING;

LABEL
:
assert
TRUE
report
"This is a string"
severity
WARNING
;

LABEL
:
assert
TRUE
report
"This is a string"
;

LABEL
:
assert
TRUE
severity
WARNING
;

LABEL : assert TRUE report "This is a string" severity WARNING;

