

use IEEE.std_logic_1164.all;

use My_Lib, otherlib.my_math_stuff.multiply;

use yetanotherlib.std_logic;

