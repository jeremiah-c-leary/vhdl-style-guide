
architecture ARCH of ENTITY is

begin

  process (one, two, three) is begin


    end process;

  process (one, two,
	   three) is
  begin

 eNd  process;
  
prOCess  (one,
	  two,
	       three) is
begIN

 end proCEss;

    Process  (one,
	  two,
	       three
       ) is
  beGIn

    end  process;

proCEss (one, two, three
	  ) is
  begin

  End process;

    process (one, two, three
	    ) is
begin

  end Process;
  a<=b;
  c<=d;

proc_name : process (one, two, three) is
  begin
  end process proc_name;

end architecture ARCH;

