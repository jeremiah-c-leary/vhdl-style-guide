
architecture RTL of FIFO is

begin


  PROC_LABEL : process 
  begin
  end process PROC_LABEL;

  -- Violations below

  PROCESS_LABEL : process 
  begin
  end process PROCESS_LABEL;

end architecture RTL;
