architecture rtl of fifo is

  signal a : std_logic; -- Comment

  -- Okay comment
  signal b : std_logic_vector;

begin

  a <= b; -- Comment 1
  c <= d; -- Comment 2
  e <= f; -- Comment 3

end architecture rtl;
