
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo IS

  end component fifo;

  component fifo Is

  end component fifo;

begin

end architecture RTL;
