
ARCHITECTURE RTL OF FIFO IS

BEGIN

END ARCHITECTURE RTL;

