
architecture RTL of FIFO is

  function func1 return integer is begin end function func1;

  FUNCTION FUNC1 return INTEGER IS BEGIN END FUNCTION FUNC1;

  procedure proc1 Is begin end procedure proc1;

begin

end architecture RTL;
