
architecture RTL of FIFO is

  function func1 return integer is begin end function func1;

  function func1 return integer is begin end function func1;

  function func1 return integer is begin end function func1;

  procedure proc1 is begin End procedure proc1;

begin

end architecture RTL;
