
architecture rtl of fifo is

begin

  procedure_call_label : postponed wr_en(a, b);

  procedure_call_label : POSTPONED wr_en(a, b);

end architecture rtl;
