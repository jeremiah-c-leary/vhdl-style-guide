
architecture RTL of FIFO is

  constant c_width : INTEGER := 16;

  constant c_depth : INTEGER := 512;

  constant c_word : INTEGER := 1024;

  constant zeros : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');

  constant zeros : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');

begin

end architecture RTL;
