
entity FIFO is

end entity;

ENTITY FIFO is

end entity;

Entity FIFO is

end entity;

