
architecture RTL of FIFO is

  type t_my_type is range -5 to 5;
  type t_my_type;

  type t_my_type is range -5 to 5;
  type t_my_type;

begin

end architecture RTL;
