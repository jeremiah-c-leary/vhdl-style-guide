
architecture rtl of e is
begin

    g_0 : if true generate
        g_1 : if true generate
            signal Sig0 : bit;
            signal Sig00 : bit;
        begin

            g_2 : for i in 0 to 0 generate

            end generate g_2;

        end generate g_1;
    end generate g_0;
end architecture rtl;

