
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo

  end component fifo;

begin

end architecture RTL;
