
architecture RTL of FIFO is

  function func1 return integer is BEGIN end function func1;

  function func1 return integer is BEGIN end function func1;

  function func1 return integer is BEGIN end function func1;

begin

end architecture RTL;
