
package pkg_fifo is

end package;

package fifo is

end package;

