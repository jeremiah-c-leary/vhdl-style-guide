
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  PROCEDURE PROC1 is BEGIN END PROCEDURE PROC1;

begin

end architecture RTL;
