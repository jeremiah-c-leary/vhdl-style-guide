
architecture RTL of FIFO is begin end architecture FIFO;

-- Violations below

architecture RTL of FIFO is begin end architecture FIFO;
library ieee;

-- Last line in the file is okay
architecture RTL of FIFO is begin end architecture FIFO;
