
generic ( );

generic (

);

generic
(
)
;
