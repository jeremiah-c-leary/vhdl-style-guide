
architecture ARCH of ENTITY is

begin

  PROC_1 : process (a, b, c) is
  begin

    case boolean_1 is

      when STATE_1 =>

        null;

      when STATE_2 =>

      null;

      when STATE_3 =>

          null;

    end case;

  end process PROC_1;


end architecture ARCH;
