
architecture RTL of FIFO is

begin

  block_label : block is begin end block block_label;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK block_label;

end architecture RTL;
