
architecture RTL of FIFO is

  function func1 return integer is begin end function f_FUNC1_F;

  FUNCTION FUNC1 RETURN INTEGER IS BEGIN END FUNCTION f_FUNC1_F;

  procedure proc1 is begin end procedure Proc1;

begin

end architecture RTL;
