
architecture rtl of fifo is

  file defaultimage : load_file_type open read_mode is load_file_name;

  file defaultimage : load_file_type open read_mode is load_file_name;

  file defaultimage : load_file_type open read_mode is load_file_name;

begin

end;
