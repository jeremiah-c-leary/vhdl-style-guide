
architecture RTL of FIFO is

  signal sig1 : STD_LOGIC;
  signal sig2 : STD_LOGIC_VECTOR(3 DOWNTO 0);

  -- Violations below

  signal sig1 : STD_LOGIC;
  signal sig2 : STD_LOGIC_VECTOR(3 downto 0);


begin

end architecture RTL;
