
library ieee;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_1164.std_logic;

library std;
    use std.env.all;

library bad_lib;
    use bad_lib.bad_pkg.bad_obj;
