
use ieee.std_logic_1164.all;

use ieee.std_logic_1164.all;
