
architecture RTL of FIFO is

begin

  block_label : block is begin end block block_label;

  BLOCK_LABEL : BLOCK IS begin END BLOCK BLOCK_LABEL;

end architecture RTL;
