
library ieee;

library ieee;

