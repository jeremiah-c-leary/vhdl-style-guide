
architecture rtl of fifo is

end architecture;
