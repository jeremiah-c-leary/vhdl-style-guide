
entity fifo is end entity;
entity e_fifo is end entity;
entity fifo_a is end entity;
entity e_fifo_a is end entity;

entity FIFO is end entity;
entity e_FIFO is end entity;
entity FIFO_a is end entity;
entity e_FIFO_a is end entity;

entity fIfo is end entity;
entity e_fIfo is end entity;
entity fIfo_a is end entity;
entity e_fIfo_a is end entity;

entity Fifo is end entity;
entity e_Fifo is end entity;
entity Fifo_a is end entity;
entity e_Fifo_a is end entity;

entity MY_FIFO is end entity;
entity e_MY_FIFO is end entity;
entity MY_FIFO_a is end entity;
entity e_MY_FIFO_a is end entity;

entity my_fifo is end entity;
entity e_my_fifo is end entity;
entity my_fifo_a is end entity;
entity e_my_fifo_a is end entity;

entity MyFifo is end entity;
entity e_MyFifo is end entity;
entity MyFifo_a is end entity;
entity e_MyFifo_a is end entity;

entity myFifo is end entity;
entity e_myFifo is end entity;
entity myFifo_a is end entity;
entity e_myFifo_a is end entity;

entity MyFIFo is end entity;
entity e_MyFIFo is end entity;
entity MyFIFo_a is end entity;
entity e_MyFIFo_a is end entity;

entity myFIFo is end entity;
entity e_myFIFo is end entity;
entity myFIFo_a is end entity;
entity e_myFIFo_a is end entity;

entity myFIfo is end entity;
entity e_myFIfo is end entity;
entity myFIfo_a is end entity;
entity e_myFIfo_a is end entity;

entity MyFifO is end entity;
entity e_MyFifO is end entity;
entity MyFifO_a is end entity;
entity e_MyFifO_a is end entity;

entity myFifO is end entity;
entity e_myFifO is end entity;
entity myFifO_a is end entity;
entity e_myFifO_a is end entity;

-- Test Pascal_Snake_Case

entity MyFifo_GreenRed_Blue is end entity;
entity e_MyFifo_GreenRed_Blue is end entity;
entity MyFifo_GreenRed_Blue_a is end entity;
entity e_MyFifo_GreenRed_Blue_a is end entity;

entity My_Fifo_Green_Red_Blue is end entity;
entity e_My_Fifo_Green_Red_Blue is end entity;
entity My_Fifo_Green_Red_Blue_a is end entity;
entity e_My_Fifo_Green_Red_Blue_a is end entity;
