
use ieee.std_logic_1164.ALL;

use ieee.std_logic_1164.ALL;

