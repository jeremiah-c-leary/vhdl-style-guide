
architecture RTL of FIFO is

  procedure average_samples;

begin

  Average_samples;

  PROC1 : process () is
  begin

     AVERAGE_SAMPLES;
     AVERAGE_SaMPLES;
     aVeRAGE_SaMPLES;

  end process;

end architecture RTL;
