
architecture RTL of FIFO is

begin


  process
  begin
  end process;

  -- Violations below

  process
    begin
  end process;

  process
begin
  end process;

end architecture RTL;
