
architecture RTL of FIFO is

  type state_machine is (IDLE, WRITE, READ, DONE);

  -- Violations below

  type state_machine is (IDLE, WRITE, READ, DONE);

begin

end architecture RTL;
