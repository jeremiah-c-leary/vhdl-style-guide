
architecture RTL of FIFO is

begin

  FOR_LABEL : for i in 0 to 7 generate
  end;
  end generate;

  -- Violations below

  FOR_LABEL : for i in 0 to 7 generate
  end;
  end generate;

  FOR_LABEL : for i in 0 to 7 generate
  end;
  end generate;

end;
