
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block is

    signal sig1   : std_logic;
    constant con1 : std_logic := '0';
    file file1    : std_logic;
    alias alias1  : subtype_indicator is name;
    alias alias1  is name;

  begin
  end block BLOCK_LABEL;

end architecture RTL;
