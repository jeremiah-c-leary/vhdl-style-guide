
entity fifo is

end entity;

entity fifo is

end entity;

entity fifo is

end entity;

entity my_fifo is

end entity;

entity my_fifo is

end entity;

entity myfifo is

end entity;

entity myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity myfifp is

end entity;

entity myfifo is

end entity;

entity e_myfifo_a is

end entity;

entity e_myfifo_a is

end entity;

entity myfifo_a is

end entity;

entity myfifo_a is

end entity;

-- Test Pascal_Snake_Case

entity myfifo_greenred_blue is end entity;

entity e_my_fifo_green is end entity;

entity my_fifo_green_a is end entity;

entity e_myfifo_greenred_blue_a is end entity;
