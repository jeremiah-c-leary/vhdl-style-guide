
library ieee;
  use ieee.numeric_std.all;
  use ieee.std_logic_1164.all;

library lib1;

library lib2;

use work.registers_pkg.all;
use work.utility_pkg.all;

architecture rtl of fifo is

begin

end architecture rtl;

library lib3;

use ieee.numeric_std.all;

entity fifo is
end entity fifo;

library lib4;

use ieee.numeric_std.all;

package fifo_pkg is
end package fifo_pkg;

library lib5;

use ieee.numeric_std.all;

package body fifo_pkg_body is
end package body fifo_pkg_body;

library lib6;

use ieee.numeric_std.all;

  use lib6.my_stuff.all;
