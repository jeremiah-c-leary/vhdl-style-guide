
architecture RTL of FIFO is

begin

  process
  begin

    for_label : for index in 4 to 23 loop

    end loop;

    for_label : for index in 4 to 23 loop

    end loop;

    for_label : for index in 4 to 23 loop

    end loop;

  end process;

end;
