
PACKAGE body fifo_pkg is

end package body fifo_pkg;

PACKAGE body fifo_pkg is

end package body fifo_pkg;

