
architecture RTL of FIFO is

begin


  LABEL_PROC : process
  begin
  end process LABEL_PROC;

  -- Violations below

  LABEL_PROCESS : process
  begin
  end process LABEL_PROCESS;

end architecture RTL;
