
CONTEXT c1;

CONTEXT c2;

CONTEXT c2;
