
library IEEE;

library IEEE;

