
library ieee;
