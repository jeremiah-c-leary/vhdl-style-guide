
context c1, c1a, c1b;

context c2, c2a, c2b;

context con3, con3a;

context lib1.c1;

context LIB1.c1;
