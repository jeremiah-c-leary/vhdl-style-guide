
entity fifo is

end entity;

entity fifo is

end entity;

entity fifo is

end entity;

entity my_fifo is

end entity;

entity my_fifo is

end entity;

entity myfifo is

end entity;

entity myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity e_myfifo is

end entity;

entity myfifp is

end entity;

entity myfifo is

end entity;

entity e_myfifo_a is

end entity;

entity e_myfifo_a is

end entity;

entity myfifo_a is

end entity;

entity myfifo_a is

end entity;

