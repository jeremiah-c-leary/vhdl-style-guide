
package fifo_pkg is

  function func_a (x : boolean) return boolean;

  function func_b (x : boolean) return boolean;

  procedure proc_a (x : boolean);

  procedure proc_b (x : boolean);

end package fifo_pkg;

package body fifo_pkg is

  function func_a (x : boolean) return integer is
  begin
  end function;

  function func_b (x : boolean) return integer is
  begin
  end function;

  function func_a (x : boolean) return integer is
  begin
  end function;

  function func_b (x : boolean) return integer is
  begin
  end function;

  procedure proc_a (x : boolean) is
  begin
  end procedure proc_a;

  procedure proc_b (x : boolean) is
  begin
  end procedure proc_b;

  procedure proc_a (x : boolean) is
  begin
  end procedure;

  procedure proc_b (x : boolean) is
  begin
  end procedure;

end package body fifo_pkg;
