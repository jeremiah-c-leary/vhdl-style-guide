
architecture RTL of FIFO is

  signal sig1 : std_logic;
  signal sig2 : std_logic;

  -- Violations below

  SIGNAL sig1 : std_logic;
  SIGNAL sig2 : std_logic;


begin

end architecture RTL;
