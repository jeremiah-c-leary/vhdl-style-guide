
library ieee;

library ieee;  --comment

-- Violations below

library ieee;

library ieee;  -- comment

library ieee;  -- comment
