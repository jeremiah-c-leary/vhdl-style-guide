
package fifo_pkg is

  attribute mark_debug of wr_en        : signal is "true";
  attribute mark_debug of almost_empty : signal is "true";
  attribute mark_debug of full         : signal is "true";

end package;
