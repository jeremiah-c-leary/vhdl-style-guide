

architecture RTL of ENTITY1 is

begin

end architecture RTL;



architecture RTL of ENTITY1 is

begin

end;


architecture RTL of ENTITY1 is

begin

end architecture;


architecture
RTL
of
ENTITY1
is
begin
end
architecture
RTL
;
