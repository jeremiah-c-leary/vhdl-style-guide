
architecture RTL OF ENT is
begin
end RTL;

architecture RTL OF ent is
begin
end rtl;

architecture RTL OF Ent is
begin
end Rtl;

architecture RTL OF ENT is
begin
end;

architecture RTL OF ENT is
begin
end architecture;

