architecture rtl of fifo is

  procedure average_samples (
    sample                 : signed;
    constant num_samples   : in integer := 0;
    file my_file           : text;
    variable sample_number : in integer;
    signal sample          : out std_logic
  );

  procedure average_samples (sample : signed; constant num_samples : in integer := 0; file my_file : text; variable sample_number : in integer; signal sample : out std_logic
 );

  procedure average_samples (
    sample : signed; constant num_samples : in integer := 0; file my_file : text; variable sample_number : in integer; signal sample : out std_logic
 );

  procedure average_samples (sample : signed; constant num_samples : in integer := 0; file my_file : text; variable sample_number : in integer; signal sample : out std_logic
  );

  procedure average_samples (
    sample                 : signed;
    constant num_samples   : in integer := 0;
    file my_file           : text;
    variable sample_number : in integer;
    signal sample          : out std_logic
 );

  procedure average_samples
  (
    sample                 : signed;
    constant num_samples   : in integer := 0;
    file my_file           : text;
    variable sample_number : in integer;
    signal sample          : out std_logic
 );

  procedure average_samples (
    sample                 : signed
    ;
    constant num_samples   : in integer := 0
;
    file my_file           : text

    ;
    variable sample_number : in integer;

    signal sample          : out std_logic
  );

begin

end architecture;
