

use IEEE.std_logic_1164.all;

use MY_LIB, OTHERLIB.my_math_stuff.multiply;

use YETANOTHERLIB.std_logic;

