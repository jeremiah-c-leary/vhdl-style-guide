
context name1;

context name2, name3;

context name4, name5, name6;

