
architecture RTL of FIFO is

begin

  process
  begin

    loop

    end loop;

    -- Violations below

    loop end loop
    ;

  end process;

end;
