
architecture RTL of FIFO is

begin

  block_label : block is BEGIN end block block_label;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
