
entity FIFO is

end entity;

entity FIFO is

end entity;

entity FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MYFIFO is

end entity;

entity MYFIFO is

end entity;

