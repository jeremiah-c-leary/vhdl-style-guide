
library ieee;

library       ieee;
