
architecture RTL of FIFO is

begin

  block_label : block IS begin end block block_label;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
