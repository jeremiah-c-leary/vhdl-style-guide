
architecture RTL of FIFO is

begin

  block_label : block is begin end block block_label;

  block_label : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
