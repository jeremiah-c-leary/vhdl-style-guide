
architecture RTL of FIFO is

  subtype counter_t is unsigned(4 downto 0);
  subtype counter is unsigned(4 downto 0);
  constant width : integer := 32;

  subtype counter is unsigned(4 downto 0);
  subtype counter_t is unsigned(4 downto 0);
  constant width : integer := 32;

begin

end architecture RTL;
