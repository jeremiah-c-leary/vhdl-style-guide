
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    null;

    NULL_LABEL : null;

  end process;

end architecture RTL;
