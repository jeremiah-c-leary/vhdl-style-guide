
architecture RTL of FIFO is

  attribute max_delay : time;

  attribute MAX_DELAY : TIME;

begin

end architecture RTL;
