
architecture rtl of fifo is

begin

  process begin

    LOOP end loop;

    LOOP END LOOP;

  end process;

end;
