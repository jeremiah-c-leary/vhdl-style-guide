
architecture RTL of FIFO is

  constant c_width : integer := 16;
  constant c_depth :   integer := 512;
  constant c_word :integer := 1024;

begin

end architecture RTL;
