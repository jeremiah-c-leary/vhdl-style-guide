
architecture rtl of fifo is

begin

  gen_test : for gv_param in t_range generate
  end generate gen_test;

  my_proc : process is
  begin

    for lv_param in t_range loop
    end loop;

  end process my_proc;

  gen_test : for GV_PARAM in t_range generate
  end generate gen_test;

  my_proc : process is
  begin

    for LV_PARAM in t_range loop
    end loop;

  end process my_proc;

end;
