package test is

  type flag_pt is PROTECTED
  end protected;

  type flag_pt is PROTECTED
  end protected;

end package test;

architecture rtl of test is

  type flag_pt is PROTECTED
  end protected;

  type flag_pt is PROTECTED
  end protected;

begin

end architecture rtl;
