
architecture rtl of fifo is

begin

  process begin

    for x in (11 downto 0) loop end loop;

    for x in (11 downto 0) loop end loop;

  end process;

end;
