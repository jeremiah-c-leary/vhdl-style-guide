
library ieee;

library IEEE;
