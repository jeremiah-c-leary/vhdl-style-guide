
package body pkg_fifo is

end package body pkg_fifo;

package body fifo is

end package body fifo;
