
architecture rtl of fifo is

  alias designator : subtype_indication is name;

  alias designator     is name;

  alias designator : subtype_indication is name;

  alias designator : (subtype_indication) is name;

begin

end architecture rtl;
