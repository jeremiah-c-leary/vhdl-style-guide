
entity fifo is

end entity;

entity fifo is

end entity;

entity fifo is

end entity;

