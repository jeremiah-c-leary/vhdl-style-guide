
architecture RTL of FIFO is

  subtype read_size is range 0 to 9;

  -- Violations below

  subtype read_size is range 0 to 9;
  subtype read_size is range 0 to 9;

begin

end architecture RTL;
