
package pack1 is new pack_name
  generic map (
    A => B,
    C => D,
    E, F
  );

package pack2 is new pack2_name;

