
use My_Math_Stuff.MY_STRING_STUFF.my_string_stuff;

use My_Math_Stuff.My_Math_Stuff.my_math_stuff;

use My_Logic_Stuff.my_logic_stuff.my_logic_stuff;

use ieee.std_logic_1164.all;
