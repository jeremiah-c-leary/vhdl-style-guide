
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block begin end block;


  BLOCK_LABEL : block begin end block;

  BLOCK_LABEL : block--Comment
    begin end block;

  BLOCK_LABEL : block --Comment
    begin end block;

  BLOCK_LABEL : block --Comment
 begin end block;

  BLOCK_LABEL : block (guard_condition)begin end block;

  BLOCK_LABEL : block (guard_condition) begin end block;

  BLOCK_LABEL : block (guard_condition)
    begin end block;

  BLOCK_LABEL : block
    begin end block;

end architecture RTL;
