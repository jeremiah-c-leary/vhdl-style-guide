
architecture rtl of fifo is

begin

  block_label : block is
  begin

  end block block_label;

------------------------------<-    80 chars    ->------------------------------
--! FPGA RX to Avalon-ST TX interface
--------------------------------------------------------------------------------

  ------------------------------<-    80 chars    ->------------------------------
  --------------------------------------------------------------------------------

  ------------------------------<-    80 chars    ->------------------------------

------------------------------<-    80 chars    ->------------------------------
--! FPGA RX to Avalon-ST TX interface
--! FPGA RX to Avalon-ST TX interface
--! FPGA RX to Avalon-ST TX interface
--------------------------------------------------------------------------------

------------------------------<-    80 chars    ->------------------------------
--! FPGA RX to Avalon-ST TX interface
--! FPGA RX to Avalon-ST TX interface
--! FPGA RX to Avalon-ST TX interface
--! FPGA RX to Avalon-ST TX interface
--------------------------------------------------------------------------------

end architecture rtl;
