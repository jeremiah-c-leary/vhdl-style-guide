
architecture RTL of FIFO is

begin

  blk_block_label : block is begin end block blk_block_label;

  block_label : block is begin end block block_label;

end architecture RTL;
