

architecture ARCH of ENTITY is

begin

end ARCH;

  architecture ARCH of ENTITY is

begin

end ARCH
architecture  ARCH  of  ENTITY  is

begin

end ARCH

  Architecture ARch Of entity Is

 begin

end ArCh

architecture ARch
 of ENTITY is

begin

end ARCH

