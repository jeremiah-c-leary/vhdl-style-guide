
architecture RTL of FIFO is

begin

  block_label : block is begin end block BLOCK_LABEL;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
