
architecture RTL of FIFO is

  procedure PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) is
   begin
   end procedure PARITY;

  procedure PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) is
   begin
   end procedure;

  procedure PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) is
   begin
   end PARITY;

  procedure PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) is
   begin
   end;

  function PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) return integer is
   begin
   end function PARITY;

  function PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) return string is
   begin
   end function;

  function PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) return natural is
   begin
   end PARITY;

  function PARITY
   (signal X : in std_logic_vector;
    signal Y : out std_logic) return positive is
   begin
   end;

begin


end architecture RTL;
