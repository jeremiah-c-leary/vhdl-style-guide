
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  procedure PROC1 IS BEGIN END PROCEDURE PROC1;

begin

end architecture RTL;
