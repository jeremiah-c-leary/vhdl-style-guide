
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    PROC_LABEL : proc(a, b, c);

    PROC_LABEL : proc;

    proc(a, b, c);

    proc;

  end process;

end architecture RTL;
