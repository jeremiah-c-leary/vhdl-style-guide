
architecture rtl of fifo is

  file defaultimage : load_file_type open read_mode is load_file_name;

  file DEFAULTIMAGE : load_file_type open read_mode is load_file_name;

  file DefaultImage : load_file_type open read_mode is load_file_name;

begin

end;
