
entity FIFO is

end entity;
architecture rtl of fifo is
begin
end architecture;

entity FIFO is
end entity;
 architecture rtl of fifo is begin end architecture;

