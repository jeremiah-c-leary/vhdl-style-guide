
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  COMPONENT fifo --Some Comemnt
  is -- Some COmment

  end component fifo;

  Component fifo--Other comment
  -- Some Comment
 is

  end component fifo;

begin

end architecture RTL;
