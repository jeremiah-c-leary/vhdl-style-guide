
architecture RTL of FIFO is

begin


  process (a, b)
  begin
  end process;

  process is
  begin
  end process;

  process begin
  end process;

  -- Violations below

  process (a, b)
  begin
  end process;

  process (a, b)
  begin
  end process;

  process is
  begin
  end process;

  process begin
  end process;

end architecture RTL;
