
architecture RTL of FIFO is

  attribute coordinate of others : COMPONENT is (0.0, 17.5);

  attribute coordinate of others : COMPONENT is (0.0, 17.5);

begin

end architecture RTL;
