
architecture rtl of fifo is

begin

  process is begin
    exit;

      exit;

  exit;

  end process;

end architecture rtl;
