
entity fifo is

begin

end entity fifo;


entity fifo is

begin

end;

entity fifo is

begin

end entity;

entity
fifo
is
begin
end
entity
fifo
;
