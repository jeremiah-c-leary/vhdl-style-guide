
configuration CFG of FIFO is

  group group1_identifier : group1_template_name ( group_constituent1 );

  group group2_identifier : group2_template_name ( group_constituent1, group_constintuent2 );

end configuration CFG;

