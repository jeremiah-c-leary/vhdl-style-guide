
architecture rtl of fifo is

  component my_block is
  end component;

  -- synthesis translate_on

  component my_block is
  end component;
  -- synthesis translate_on

begin

end architecture;
