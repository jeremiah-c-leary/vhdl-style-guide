
architecture RTL of FIFO is

  attribute MAX_DELAY : time;

  ATTRIBUTE MAX_DELAY : TIME;

begin

end architecture RTL;
