
architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end;

