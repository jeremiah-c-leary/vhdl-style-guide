
architecture rtl of fifo is

begin

  process begin

    loop END loop;

    LOOP END LOOP;

  end process;

end;
