
architecture RTL of ENT is
begin
end architecture RTL;

architecture RTL of ENT is
begin
end rtl;

architecture RTL of ENT is
begin
end architecture Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;

