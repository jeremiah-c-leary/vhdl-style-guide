
------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

architecture rtl of fifo is

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

begin

  process

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

  begin

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

  end process;

end architecture rtl;

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

