
architecture rtl of fifo is

begin

  process begin

    WHILE condition loop end loop;

    WHILE condition loop end loop;

  end process;

end;
