
-- failure
  -- passed

architecture RTL of FIFO is

-- failure
  -- passed
    -- failure

begin

-- failure
  -- passed
    -- failure

end architecture RTL;
