
entity FIFO is

end entity;


entity FIFO is

end entity;


entity FIFO2 is

end entity ;
