
architecture RTL of ENT is begin end architecture RTL;

architecture RTL of

ENT is
begin
end;

architecture RTL of
-- Some domment
 ENT is
begin
end;

architecture RTL of--some comment
 ENT is
begin
end;

