architecture ARCH of FIFO is

  signal sig1 : std_logic;        -- comment
  signal sig1 : std_logic;    -- comment
  signal sig1 : std_logic;  -- comment
  signal sig1 : std_logic;         -- comment
  signal sig1 : std_logic; -- comment
  -- This comment should be left alone
  signal sig1 : std_logic;     -- comment
  signal sig1 : std_logic;     -- comment
  signal sig1 : std_logic; -- comment
  signal sig1 : std_logic;            -- comment
  signal sig1 : std_logic;    -- comment

  signal sig1 : std_logic;      -- comment
  signal sig1 : std_logic;     -- comment
  signal sig1 : std_logic; -- comment
  signal sig1 : std_logic;       -- comment
  signal sig1 : std_logic;   -- comment
  -- This comment should be left alone
  signal sig1 : std_logic;      -- comment
  signal sig1 : std_logic;     -- comment
  signal sig1 : std_logic; -- comment
  signal sig1 : std_logic;            -- comment
  signal sig1 : std_logic;   -- comment

  --------------------
  -- COMMENT BLOCK
  --
  --
  --
  --------------------

begin

end architecture ARCH;
