
architecture rtl of fifo is

  procedure proc is
  begin
  end proc;

  procedure proc is
  begin
  end proc;

  function func return integer is
  begin
  end func;

  function func return integer is
  begin
  end;

  procedure proc;

  function func return integer is
  begin
  end;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end proc;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end proc;

begin

end architecture rtl;
