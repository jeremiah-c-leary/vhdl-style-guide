
architecture rtl of fifo is

  alias a_designator is name;

  alias designator is name;

begin

end architecture rtl;
