
package body fifo_pkg is

end package body;

package  body fifo_pkg is

end package body;

package body fifo_pkg  is

end package body;

package  body  fifo_pkg  is

end package body;
