
entity ENTITY1 is
  port (
    PORT1 : in    std_logic;
    PORT2 : out   std_logic;
    PORT3 : inout std_logic;
    PORT4 : in    std_logic;
    PORT5 : out   std_logic;
    PORT6 : inout std_logic
  );
end entity ENTITY1

architecture ARCH of ENTITY1 is

begin

end architecture ARCH;
