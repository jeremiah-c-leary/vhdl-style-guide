
attribute LOCATION: COORDINATE;

attribute PIN_NO: POSITIVE;

