
architecture RTL of FIFO is

  function func1 (
    a : integer;
    b: integer
  ) return integer;

  function func1 (
a : integer;
    b: integer
  ) return integer;

  function func1 (a : integer;b: integer) return integer;

begin

end architecture RTL;
