
architecture RTL of FIFO is

shared variable Counter: SharedCounter;

shared variable addend, augend, result: ComplexNumber := "asdf";

shared
variable
addend
,
augend
,
result
:
ComplexNumber
;

begin

end architecture RTL;
