
architecture RTL of ENT IS
begin
end RTL;

architecture RTL of ent IS
begin
end rtl;

architecture RTL of Ent IS
begin
end Rtl;

architecture RTL of ENT IS
begin
end;

architecture RTL of ENT IS
begin
end architecture;

