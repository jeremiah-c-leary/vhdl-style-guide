
--------------------------------------------------------------------------------
-- Comment
-- Comment
-- Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--+ Comment
--+ Comment
--+ Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--| Comment
--| Comment
--| Comment
--| Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--!-- Comment
--!-- Comment
--!-- Comment
--!-- Comment
--------------------------------------------------------------------------------

-- comment
-- comment
