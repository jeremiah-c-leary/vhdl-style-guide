
architecture RTL of FIFO is

  attribute max_delay : time;

  ATTRIBUTE max_delay : TIME;

begin

end architecture RTL;
