
package body fifo is

end package body fifo;

package body fifo is

end;

package body fifo is

end package body;

package
body
fifo
is
end
package
body
fifo
;
