--
-- This should pass
--| This should pass
----------This should pass
--==================

-- This should fail
--| This should fail
----------This should pass
--
--==================


--¨

