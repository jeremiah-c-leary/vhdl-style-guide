
library ieee;

  library ieee;
