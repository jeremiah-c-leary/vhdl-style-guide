
architecture rtl of fifo is

begin

  test1 <= 1 after 10 ns;

  test1 <= 1 after 10 ns;

end architecture;
