
architecture RTL of FIFO is

  function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

  pure function func1 (a : integer) return integer is
  begin
  end;

  impure function func1 (a : integer) return integer is
  begin
  end;

  -- Fixes follow

  function func1 return integer is
  begin
  end;

  function func1 return integer is
  begin
  end;

  function func1 return integer is
  begin
  end;

  function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  pure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  impure function func1 return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

  function func1 (a : integer) return integer is
  begin
  end;

begin

end architecture RTL;
