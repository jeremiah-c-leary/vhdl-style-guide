
architecture RTL of FIFO is

  subtype counter is unsigned(4 downto 0);

  -- Violations below

  subtype counter    is unsigned(4 downto 0);

begin

end architecture RTL;
