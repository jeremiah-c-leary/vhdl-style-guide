
architecture RTL of FIFO is

  signal sig1,                sig2 : std_logic;
  signal sig2,                sig3 : std_logic;



  signal signal1a,            signal1b : std_logic;
  signal sig2a,               sig2b : std_logic;
  -- Comment line separating signals
  signal really_long_name,    shorter_name : std_logic;
  signal short_name,          some_other_really_long_name: std_logic;

  -- Blank line separating signals

  signal name,                name2 : std_logic;

  signal very_very_long_name, some_other name : std_logic;
  signal short_name2,         short_name3 : std_logic;

begin

end architecture RTL;
