
architecture RTL of FIFO is





  alias ident : std_logic_vector(3 downto 0) is write_enable [name1, name2 return integer];

  alias ident : std_logic_vector(3 downto 0) is write_enable [name1, name2];

  alias ident : std_logic_vector(3 downto 0) is write_enable [return integer];

  alias ident : std_logic_vector(3 downto 0) is write_enable;


  alias ident is write_enable [name1, name2 return integer];

  alias ident is write_enable [name1, name2];

  alias ident is write_enable [return integer];

  alias ident is write_enable;

begin

end architecture RTL;
