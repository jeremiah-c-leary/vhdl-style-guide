
entity FIFO is

end entity;

entity FIFO IS

end entity;

entity FIFO Is

end entity;
