
architecture RTL of FIFO is

  function func_1 ()

begin

  OUT1 <= Func_1;

  PROC1 : process () is
  begin

     sig1 <= FUNC_1;

  end process;

end architecture RTL;

