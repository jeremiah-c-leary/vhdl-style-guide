
architecture rtl of fifo is

begin

  x <= a sll b srl c sla d sra e rol f ror g;

  x <= a sll b srl c sla d sra e rol f ror g;

end architecture;
