
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--+-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|---------------------------------[ abcdef ]==================================

--------------------------------------------------------------------------------
-- Comment
--|-[ abcdef ]==================================================================

--------------------------------------------------------------------------------
-- Comment
--|------------------------------------------------------------------[ abcdef ]=

  ------------------------------------------------------------------------------
  -- Comment
  --+---------------------------------------------------------------------------

-- comment
-- comment

--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
