

use ieee.std_logic.1164;

use ieee.std_logic.1164, ieee.std_logic_arith.all;

use ieee.std_logic."ceil";

use ieee.std_logic."ceil", ieee.std_logic."ceil";
