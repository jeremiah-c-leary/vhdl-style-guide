
architecture RTL of FIFO is

  signal sig1 : std_logic;

  -- Violations below

  signal sig1 : std_logic := '1';


begin

end architecture RTL;
