
architecture RTL of FIFO is

  attribute max_delay : time;
  attribute max_delay     : time;

  -- Violations below

  attribute max_delay: time;

begin

end architecture RTL;
