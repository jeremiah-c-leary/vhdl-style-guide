
entity fifo is

end;

architecture rtl of fifo is
begin
end;
