
entity FIFO is

end entity FIFO;


entity FIFO is

end entity;


entity FIFO2 is

end entity ;
