
architecture RTL of FIFO is

  type state_machine_t is (idle, write, read, done);
  type state_machine is (idle, write, read, done);

  constant width : integer := 32;

  type state_machine_t is (idle, write, read, done);
  type state_machine;

  constant width : integer := 32;

  type state_machine is (idle, write, read, done);
  type state_machine_t is (idle, write, read, done);

  constant width : integer := 32;

  type state_machine;
  type state_machine_t is (idle, write, read, done);

  constant width : integer := 32;

begin

end architecture RTL;
