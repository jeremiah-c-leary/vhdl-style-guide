
architecture RTL of FIFO is

  variable   c_width : integer := 16;
  variable c_depth : integer := 512;
  variable     c_word : integer := (12, 13, 15);

begin

  process

    variable   c_width : integer := 16;
    variable c_depth : integer := 512;
    variable  c_word : integer := (12, 13, 15);
    variable          c_word : integer := (12, 13, 15);

  begin end process;

end architecture RTL;
