
architecture RTL of FIFO is

  procedure proc1 is begin end procedure PROC1;

  PROCEDURE PROC1 IS BEGIN END PROCEDURE PROC1;

  function func1 return integer is begin end function Func1;

begin

end architecture RTL;
