
package pkg_fifo is

end package pkg_fifo;

package fifo is

end package fifo;
