
entity fifo is

end entity;

entity FIFO is

end entity;

entity Fifo is

end entity;

