
architecture RTL of FIFO is

  function func1 return integer is begin end function F_func1_f;

  FUNCTION FUNC1 RETURN INTEGER IS BEGIN END FUNCTION F_func1_f;

  procedure proc1 is begin end procedure Proc1;

begin

end architecture RTL;
