
--This should pass
context CON1 is

end context CON1;

--These should fail
context CON1 is
end context con1;

context CO1 is

end context Con1;
