
architecture rtl of fifo is

begin

  process is begin
    exit;

    exit;

    exit_label : exit;

    exit_label : exit;

  end process;

end architecture rtl;
