
architecture rtl of fifo is begin end architecture rtl;

architecture rtl of fifo is begin end architecture rtl;

architecture rtl    of fifo is begin end architecture rtl;

architecture rtl of    fifo is begin end architecture rtl;

architecture rtl of fifo    is begin end architecture rtl;

