
use My_Math_Stuff.my_string_stuff.my_math_stuff;

use My_Math_Stuff.my_math_stuff.my_math_stuff;

use My_Logic_Stuff.my_logic_stuff.MY_MATH_STUFF;
