
architecture arch of entity1 is

begin

  block_label : block is
  
    type type1 is access subtype_indication more other;

  begin
  
  end block block_label;

end architecture arch;
