
architecture RTL of FIFO is

  procedure proc1 is begin END procedure proc1;

  PROCEDURE PROC1 IS BEGIN END PROCEDURE PROC1;

begin

end architecture RTL;
