
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--+-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|--------------------------------[ abcdef ]===================================

--------------------------------------------------------------------------------
-- Comment
--|-[ abcdef ]==================================================================

--------------------------------------------------------------------------------
-- Comment
--|------------------------------------------------------------------[ abcdef ]=

architecture rtl of fifo is

  ------------------------------------------------------------------------------
  -- Comment
  --+---------------------------------------------------------------------------

begin

end architecture rtl;

-- comment
-- comment

--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
