

architecture ARCH of ENTITY1 is

begin

end architecture;
