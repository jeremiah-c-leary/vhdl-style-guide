--
-- This should pass
--| This should pass
----------This should pass
--==================

--This should fail
--|This should fail
----------This should pass
--
--==================


--¨

-- pragmas should be ignored
--vhdl_comp_off
--vhdl_comp_on

