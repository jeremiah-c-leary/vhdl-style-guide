
architecture RTL of FIFO is

  procedure proc1 is
  begin
  end procedure proc1;

  procedure proc1 is
  begin
  end procedure;

  procedure proc1 is
  begin
  end proc1;

  procedure proc1 is
  begin
  end;

  -- Fixes follow

  procedure proc1 is
  begin
  end     procedure proc1;

  procedure proc1 is
  begin
  end procedure      proc1;

  procedure proc1 is
  begin
  end     procedure      proc1;

  procedure proc1 is
  begin
  end     procedure;

  procedure proc1 is
  begin
  end     proc1;

begin

end architecture RTL;
