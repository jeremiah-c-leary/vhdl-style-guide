
architecture RTL of FIFO is

  signal sig1 : std_logic_vector(3 downto 0);
  constant c_cons1 : integer := 200;
  constant c_cons2 : integer := 200;

begin


end architecture RTL;

