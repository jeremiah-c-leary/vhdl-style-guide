
architecture RTl of FIFO is

  component fifo is

  end component;

  component fifo is

  end component;

begin

end architecture RTL;
