
architecture rtl of fifo is

  alias designator is name;

  ALIAS designator is name;

begin

end architecture rtl;
