
architecture RTL of FIFO is

begin

  PROC_LABEL : postponed process is
  begin

  end process PROC_LABEL;

  PROC_LABEL : postponed process is
  begin

  end process PROC_LABEL;

  PROC_LABEL : postponed process is
  begin

  end process PROC_LABEL;

  PROC_LABEL : process is
  begin

  end process PROC_LABEL;

  PROC_LABEL : process is
  begin

  end process PROC_LABEL;

end architecture RTL;
