
architecture rtl of fifo is

begin

  process begin

    for x IN (31 downto 0) loop end loop;

    for x IN (31 downto 0) loop end loop;

  end process;

end;
