
package fifo_pkg is

end package fifo_pkg;

package fifo_pkg is

end package fifo_pkg;

package fifo_pkg is

end fifo_pkg;

