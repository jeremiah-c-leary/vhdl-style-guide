
library ieee;

library fifo, ram;

library gates;


library ieee;
 library fifo, ram;
 library gates;
