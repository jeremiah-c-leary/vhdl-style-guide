
architecture RTL of FIFO is

  function func1 return integer is begin

    loop

      NULL;
      null_label : NULL;

    end loop;

  end function func1;

  function func1 return integer is begin

    loop

      NULL;
      null_label : NULL;

    end loop;

  end function func1;

begin

end architecture RTL;
