
architecture RTL of FIFO is

  CONSTANT c_width : integer := 16;

  CONSTANT c_depth : integer := 512;

  CONSTANT c_word : integer := 1024;

begin

end architecture RTL;
