
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate
    -- Comment
    when choice =>
      -- Comment
      a <= 0;

    -- Comment
    when choice =>
      -- Comment
      a <= 0;

      -- Comment

  end generate;

  GEN_LABEL : case expression generate
-- Comment
    when choice =>
         -- Comment
      a <= 0;

       -- Comment
    when choice =>
   -- Comment
      a <= 0;

  -- Comment

  end generate;


end architecture;
