
library     ieee;
