
architecture rtl of fifo is

begin

  process begin

    loop end LOOP;

    LOOP END LOOP;

  end process;

end;
