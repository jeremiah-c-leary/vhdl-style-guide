
context c1;

context    c2;

context my_lib.c1;

context    my_lib.c2;
