
use stdio.all;

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.std_logic_arith.all;


library ieee;
  use ieee.std_logic_1164.all;
use work.registers_pkg.all;
use work.utility_pkg.all;

-- Entity declaration

entity fifo is end;
use work.utility_pkg.all;

entity fifo is end;
use work.utility_pkg.all;

-- context

context selected_name;
use work.utility_pkg.all;

context selected_name;
use work.utility_pkg.all;

-- package declaration

package fifo_pkg is end package;
use work.utility_pkg.all;

package fifo_pkg is end package;
use work.utility_pkg.all;

-- configuration

configuration fifo_cfg of fifo is end configuration;
use work.utility_pkg.all;

configuration fifo_cfg of fifo is end configuration;
use work.utility_pkg.all;

-- package

package fifo_pkg is new fifo_pkg;
use work.utility_pkg.all;

package fifo_pkg is new fifo_pkg;
use work.utility_pkg.all;

-- context declaration

context my_context is end;
use work.utility_pkg.all;

context my_context is end;
use work.utility_pkg.all;

-- architecture

architecture rtl of fifo is begin end;
use work.utility_pkg.all;

architecture rtl of fifo is begin end;
use work.utility_pkg.all;

-- package body

package body fifo_pkg is end package body;
use work.utility_pkg.all;

package body fifo_pkg is end package body;
use work.utility_pkg.all;

