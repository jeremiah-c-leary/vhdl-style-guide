
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo

  end component fifo;

  component
    fifo

  end component fifo;

  component fifo--Comment
  end component fifo;

  component fifo--Comment
   is end component fifo;

begin

end architecture RTL;
