
architecture RTL of FIFO is

begin


  PROCESS
  begin
  end process;

  -- Violations below

  PROCESS
  begin
  end process;

end architecture RTL;
