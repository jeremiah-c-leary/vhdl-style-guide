
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate
    when choice =>

  end generate;

  GEN_LABEL : case expression generate
    when choice =>

  end generate;

end architecture;
