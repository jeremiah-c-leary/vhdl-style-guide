
entity FIFO is
  port (
    I_INPUT : in std_logic
  );
end entity FIFO;


entity FIFO is
  port (
    I_INPUT : in std_logic
  );
 end entity FIFO;

entity FIFO is
  port (
    I_INPUT : in std_logic
  );
end entity FIFO;
