library ieee;

package body fifo_pkg is

end package body;

-- Violation below

package body fifo_pkg is

-- Comments are not allowed

end package body;


library ieee;
package body fifo_pkg is

  constant a : std_logic;

end package body;

