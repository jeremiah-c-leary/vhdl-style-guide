
architecture RTL of ENT is
begin
end RTL;

architecture RTL of ent is
begin
end rtl;

architecture RTL of Ent is
begin
end Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;

