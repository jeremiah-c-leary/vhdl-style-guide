
--------------------------------------------------------------------------------
-- Comment
-- Comment
-- Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--+ Comment
--+ Comment
--+ Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--| Comment
--| Comment
--| Comment
--| Comment
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--!-- Comment
--!-- Comment
--!-- Comment
--!-- Comment
--------------------------------------------------------------------------------

-- comment
-- comment
-- comment
-- comment
-- comment


--+ Comment
--+ Comment
--+ Comment


--| Comment
--| Comment
--| Comment
--| Comment

  ------------------------------------------------------------------------------
  --+ Comment
  --+ Comment
  --+ Comment
  ------------------------------------------------------------------------------
