
architecture RTL of ENTITY1 is

  subtype range_st is integer range 0 to 9;
  subtype width_st is integer range 16 to 128;

  subtype range_subt is integer range 0 to 9;
  subtype width_subt is integer range 16 to 128;

  subtype rangest is integer range 0 to 9;
  subtype widthst is integer range 16 to 128;

begin

end architecture RTL;
