
architecture RTL of FIFO is

begin

  block_label : block is begin end block block_label;

  BLOCK_LABEL : BLOCK is BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
