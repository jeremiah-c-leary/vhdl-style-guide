

architecture ARCH of ENTITY is

  signal e_sig1, d_sig2 : std_logic;
  signal a_sig10, c_sig2 : std_logic;
  signal b_sig100, b_sig2 : std_logic_vector (31 downto 0);
  signal c_sig1000, a_sig2 : std_logic;
  
  signal e_sig100,    d_sig2 : std_logic;
  signal a_sig1000,   c_sig2 : std_logic;
  signal b_sig10000,  b_sig2 : std_logic_vector (31 downto 0);
  signal c_sig100000, a_sig2 : std_logic;

begin

end architecture ARCH;

architecture ARCH of ENTITY is

  signal e_sig12,      d_sig2 : std_logic;
  signal a_sig120,     c_sig2 : std_logic;
  signal b_sig1200,    b_sig2 : std_logic_vector (31 downto 0);
  signal c_sig12000,   a_sig2 : std_logic;
  
  signal e_sig1200,    d_sig2 : std_logic;
  signal a_sig12000,   c_sig2 : std_logic;
  signal b_sig120000,  b_sig2 : std_logic_vector (31 downto 0);
  signal c_sig1200000, a_sig2 : std_logic;

  signal a, b ,c : std_logic;

begin

end architecture ARCH;
