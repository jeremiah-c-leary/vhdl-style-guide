
architecture RTL of FIFO is

  constant c_width : integer := 16;

  constant C_DEPTH : integer := 512;

  constant C_word : integer := 1024;

begin

end architecture RTL;
