
architecture RTL of FIFO is

  ATTRIBUTE ram_init_file : string;
  ATTRIBUTE ram_init_file of ram_block :
    signal is "contents.mif";

  ATTRIBUTE ram_init_file : string;
  ATTRIBUTE ram_init_file of ram_block :
    signal is "contents.mif";

  ATTRIBUTE ram_init_file : string;
  ATTRIBUTE ram_init_file of ram_block :
    signal is "contents.mif";

begin

end architecture RTL;
