
architecture rtl of fifo is

  alias DESIGNATOR is name;

  alias DESIGNATOR is name;

begin

end architecture rtl;
