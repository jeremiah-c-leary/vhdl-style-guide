

entity FIFO is
  port (
    port1 : in std_logic;
    port1 : out std_logic;
    port1 : inout std_logic bus;
    port1 : buffer std_logic bus := "asdf";
    port1 : linkage std_logic := "asdf";
    port1 : std_logic
  );
end entity FIFO;

entity FIFO is
  port (
    signal port1 : in std_logic;
    signal port1 : out std_logic;
    signal port1 : inout std_logic;
    signal port1 : buffer std_logic;
    signal port1 : linkage std_logic;
    signal port1 : std_logic
  );
end entity FIFO;
