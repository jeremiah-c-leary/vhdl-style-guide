
entity FIFO IS

end entity;

entity FIFO IS

end entity;

entity FIFO IS

end entity;

