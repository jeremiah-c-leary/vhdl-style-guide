
architecture RTL of FIFO is

begin

  IF_LABEL : if a = '1' GENERATE

  elsif b = '1' GENERATE

  else GENERATE

  end generate;

  -- Violations below

  IF_LABEL : if a = '1' GENERATE

  elsif b = '1' GENERATE

  else GENERATE

  end generate;

end;
