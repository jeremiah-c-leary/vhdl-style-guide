
package body test is

  type flag_pt is protected body
  end PROTECTED body;

  type flag_pt is protected body
  end PROTECTED body;

end package body test;

architecture rtl of test is

  type flag_pt is protected body
  end PROTECTED body;

  type flag_pt is protected body
  end PROTECTED body;

begin

end architecture rtl;
