
architecture rtl of fifo is

  file defaultImage : load_file_type open read_mode is load_file_name;

  file defaultImage : load_file_type open read_mode is       load_file_name;

begin

end architecture rtl;
