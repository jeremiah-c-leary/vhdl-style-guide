
architecture rtl of fifo is

begin

  process begin

    report "hello" SEVERITY FAILURE;

    report "hello" severity FAILURE;

  end process;

end architecture rtl;
