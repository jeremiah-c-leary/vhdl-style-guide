
ARCHITECTURE rtl of fifo is

begin

END RTL;
