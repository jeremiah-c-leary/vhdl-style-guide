
architecture RTL of FIFO is

begin

  block_label : block is begin end BLOCK block_label;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
