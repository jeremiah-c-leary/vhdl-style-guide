
architecture RTL of FIFO is

  function func1 return integer is begin end function func1;

  FUNCTION FUNC1 RETURN INTEGER IS BEGIN END FUNCTION FUNC1;

  procedure proc1 is begin end procedure Proc1;

begin

end architecture RTL;
