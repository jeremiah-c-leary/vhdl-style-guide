
architecture RTL of FIFO is

  signal sig1 : std_logic;

  subtype counter is unsigned(4 downto 0);

  -- Violations below

  signal sig1 : std_logic;
  subtype counter is unsigned(4 downto 0);

begin

end architecture RTL;
