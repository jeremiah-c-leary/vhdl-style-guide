
architecture ARCH of ENTITY is

  sig1        -- comment
  sig1     -- comment
  sig1   -- comment
  sig1          -- comment
  sig1  -- comment

begin

end architecture ARCH;
