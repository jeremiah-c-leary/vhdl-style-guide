
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block is
  begin
  end block;

  a <= b;

  BLOCK_LABEL : block is
  begin
  end block;

  a <= b;

end architecture RTL;
