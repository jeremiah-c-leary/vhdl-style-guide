
package fifo_pkg IS

end package;

package fifo_pkg IS

end package;

