-------------------------------------------------------------------------------
--  Next line is a failure 
--                                                                                                                        This is a failure
-------------------------------------------------------------------------------

-- Line below is a failure because the **is** is to far too the right
architecture RTL of ENT                                                                                                  is

  signal a, b, c, d, e, f, g, asf,   asfd  ,   a  , f  ,   a,  f,  e  ,e  ,f  ,a ,e  ,f , e, k, l,      f456h, a,  34pll, drt : std_logic;

signal a : std_logic_vector(15 downto 0);

begin

end architecture RTL;
