
architecture rtl of fifo is

begin

  proc_label :
  postponed
  process is
  begin
  end process;

  proc_label
  :
  postponed
  process is
  begin
  end process;

  proc_label : postponed
  process is
  begin
  end process;

  proc_label :
  process is
  begin
  end process;

  proc_label
  : process is
  begin
  end process;



end architecture rtl;
