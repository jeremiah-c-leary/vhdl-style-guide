
package BODY fifo_pkg is

end package body fifo_pkg;

package BODY fifo_pkg is

end package body fifo_pkg;

