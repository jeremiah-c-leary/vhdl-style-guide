
architecture RTL of FIFO is

begin


  process IS
  begin
  end process;

  -- Violations below

  process IS
  begin
  end process;

end architecture RTL;
