
architecture RTL of FIFO is

  signal a, b, c, d : std_logic;

  signal a, b, c, d : std_logic;

begin

  process (a, b, c, d) is
  begin
  end process;

  process (a, b, c, d) is
  begin
  end process;

  process (a,     b,    c,     d) is
  begin
  end process;

  process (a, b, c
           d, e, f) is
  begin end process;

end architecture RTL;
