
entity FIFO is

end entity fifo;

entity FIFO is

end ENTITY FIFO;

entity FIFO is

end Entity FIFO;

