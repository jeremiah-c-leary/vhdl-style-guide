
architecture RTL of FIFO is

  shared variable shar_var1 : integer;

begin

  process
    variable var1 : integer;
  begin
  end process; 

end architecture RTL;

-- Violations below

architecture RTL of FIFO is

  shared variable shar_var1 : integer := 0;

begin

  process
    variable var1 : integer := 20;
  begin
  end process; 

end architecture RTL;
