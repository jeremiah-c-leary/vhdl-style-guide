
context c1;

context    c2;

