
architecture rtl of fifo is

BEGIN

end architecture rtl;

