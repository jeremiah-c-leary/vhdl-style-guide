architecture rtl of fifo is

  alias ident is << CONSTANT dut.test : std_logic >>;
  alias ident is << CONSTANT dut.test : std_logic >>;
  alias ident is << CONSTANT dut.test : std_logic >>;

  alias ident is << signal dut.test : std_logic >>;
  alias ident is << SIGNAL dut.test : std_logic >>;
  alias ident is << Signal dut.test : std_logic >>;

  alias ident is << variable dut.test : std_logic >>;
  alias ident is << VARIABLE dut.test : std_logic >>;
  alias ident is << Variable dut.test : std_logic >>;

begin

end architecture rtl;
