
architecture RTL of FIFO is

  function func1 return integer is begin

    loop

      next_label : next my_loop when condition;
      next_label : next my_loop when condition;

    end loop;

  end function func1;

  function func1 return integer is begin

    loop

      next_label : next my_loop when condition;
      next_label : next my_loop when condition;

    end loop;

  end function func1;

begin

end architecture RTL;
