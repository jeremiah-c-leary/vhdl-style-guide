
architecture rtl of fifo is

begin

  gen_label : for X in range (3 downto 0) generate

  end generate;

  gen_label : for X in range (3 downto 0) generate

  end generate;

end architecture;
