
architecture RTL of ENT is

begin

  process
  begin

    a <= '1';
    b <= '0';

  end process;

end architecture RTL;
