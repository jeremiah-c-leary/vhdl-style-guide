
package fifo_pkg is

  signal wr_en        : std_logic; -- Comment
  signal rd_en        : std_logic; -- Comment
  constant c_constant : integer;   -- Comment

  signal wr_en : std_logic; -- Comment
  signal rd_en   : std_logic;  -- Comment
  constant c_constant : integer;         -- Comment

end package;

