
package body fifo_pkg is

end fifo_pkg;

package body fifo_pkg is

end fifo_pkg;

package body fifo_pkg is

end;

