
architecture rtl of fifo is

  procedure proc is
  begin
  end procedure proc;

  procedure proc is
  begin
  end proc;

  function func return integer is
  begin
  end function func;

  function func return integer is
  begin
  end func;

  function func return integer;

  procedure proc is
  begin
  end procedure proc;

begin

end architecture rtl;
