
architecture RTL of FIFO is

  attribute max_delay : TIME;

  ATTRIBUTE MAX_DELAY : TIME;

begin

end architecture RTL;
