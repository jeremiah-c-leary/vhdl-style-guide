
architecture RTL of FIFO is

  function func1 (a : integer) return integer;

  -- Violations follow

  function func1 (a : integer) return integer;

  function func1 (a : integer) return integer;

begin

end architecture RTL;
