
ARCHITECTURE rtl of fifo is

begin

END architecture rtl;
