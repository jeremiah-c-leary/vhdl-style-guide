
architecture RTL of ENT is
begin
end architecture RTL;

architecture RTL of ENT is
begin
end RTL;

architecture RTL of ENT is
begin
end      architecture RTL;

architecture RTL of ENT is
begin
end
architecture RTL;

