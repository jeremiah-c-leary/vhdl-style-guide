
architecture RTL of ENT is
begin
end ARCHITECTURE RTL;

architecture RTL of ENT is
begin
end rtl;

architecture RTL of ENT is
begin
end architecture Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end Architecture;
