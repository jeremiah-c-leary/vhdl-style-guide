
architecture RTL of FIFO is

  signal c_width : integer :=     16;
  signal c_depth : integer := 512;
  signal c_word : integer :=(12, 13, 15);

begin

end architecture RTL;
