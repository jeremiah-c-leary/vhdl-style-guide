
architecture rtl of fifo is

begin

  PROC_LABEL : process begin end process;

  PROC_LABEL : postponed process begin end process;

  PROC_LABEL -- Comment
  : process begin end process;

  PROC_LABEL -- Comment
  : postponed process begin end process;

  PROC_LABEL -- Comment




  : process begin end process;

  PROC_LABEL -- Comment




  : postponed process begin end process;

end;
