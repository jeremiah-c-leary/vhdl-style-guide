
architecture RTL of FIFO is

begin

  process
  begin

    FOR_LABEL : for index in 4 to 23 loop

    end loop;

    FOR_LABEL :for index in 4 to 23 loop

    end loop;

    For_label :    for index in 4 to 23 loop

    end loop;

  end process;

end;
