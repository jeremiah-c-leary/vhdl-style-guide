architecture RTL of FIFO is

  attribute LOCATION: COORDINATE;

  attribute PIN_NO: POSITIVE;

begin

end architecture RTL;
