
architecture RTL of FIFO is





  alias ident : std_logic is write_enable signature1;

  alias ident is write_enable signature1;

  alias ident : std_logic is write_enable;

  alias ident is write_enable;

  alias 'a' is write_enable;

  alias "abc" is write_enable;



begin

end architecture RTL;
