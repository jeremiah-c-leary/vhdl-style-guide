
architecture RTL of FIFO is

  SUBTYPE state_machine is subtype_indication;

  -- Violations below

  SUBTYPE state_machine is subtype_indication;

begin

end architecture RTL;
