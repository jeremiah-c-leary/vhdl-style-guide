
architecture RTL of FIFO is

  FUNCTION func1 return integer is begin end function func1;

  FUNCTION func1 return integer is begin end function func1;

  FUNCTION func1 return integer is begin end function func1;

begin

end architecture RTL;
