

context c1;

library ieee;
  context c2;

context con1 is

  library ieee;
    context c3;
end context con1;

