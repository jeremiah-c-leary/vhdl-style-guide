
use My_Math_Stuff.MY_STRING_STUFF.MY_STRING_STUFF;

use My_Math_Stuff.My_Math_Stuff.MY_MATH_STUFF;

use My_Logic_Stuff.my_logic_stuff.MY_LOGIC_STUFF;

use ieee.std_logic_1164.all;
