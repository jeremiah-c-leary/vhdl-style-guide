

architecture Arch of ENTITY is

begin

End  architecture ARCH;

  architecture ARCH of EntITY is

begin

end Architecture
architecture  ARCH  of  ENTITY  is

begin

end  architecture ARCH

 Architecture ARch Of entity Is

 begin

 eND architecture ArCh

architecture ARch
 of ENTITY is

begin

 end archITecture   ARCH

architecture ARCH of ENTITY is
begin
end architecture ARCH;

architecture ARCH of ENTITY is

begin

  process () is
  begin
  end process;

end architecture ARCH;

