
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  PROCEDURE PROC1 is BEGIN END PROCEDURE PROC1;

  FUNCTION FUNC1 RETURN INTEGER Is BEGIN END FUNCTION FUNC1;

begin

end architecture RTL;
