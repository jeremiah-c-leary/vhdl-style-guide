
architecture RTL of ENT is
BEGIN
end RTL;

architecture RTL of ENT is
begin
end rtl;

architecture RTL of ENT is
Begin
end Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;

