
package body fifo_pkg is

end PACKAGE body fifo_pkg;

package body fifo_pkg is

end PACKAGE body fifo_pkg;
