
package my_pkg IS new my_generic_pkg
  generic map (
    g_my_generic => 2
  );

package my_pkg IS new my_generic_pkg
  generic map (
    g_my_generic => 2
  );
