
architecture RTL of FIFO is

  attribute coordinate of ALL : component is (0.0, 17.5);

  attribute coordinate of ALL :component is (0.0, 17.5);

begin

end architecture RTL;
