
architecture RTL of FIFO is

begin

  process
  begin

    loop end loop LOOP_LABEL;

    LOOP_LABEL : loop end loop LOOP_LABEL;

    loop end loop;

    LOOP_LABEL1 : loop end loop LOOP_LABEL1;

  end process;

end;
