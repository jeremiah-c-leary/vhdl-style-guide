
package body fifo_pkg is

END package body fifo_pkg;

package body fifo_pkg is

END package body fifo_pkg;

