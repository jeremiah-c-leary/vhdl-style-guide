
architecture RTL of FIFO is

  type my_array is array(natural range 0 to 7) of        std_logic_vector(7 downto 0);
  type my_array is array(natural range 0 to 7) of std_logic_vector(7 downto 0);

  type my_array is array(0 to 7) of        std_logic_vector(7 downto 0);
  type my_array is array(0 to 7) of std_logic_vector(7 downto 0);

begin

end architecture RTL;
