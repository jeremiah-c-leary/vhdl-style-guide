
package fifo_pkg is

end package;

package fifo_pkg --comment
is

end package;

