
architecture RTL of FIFO is

begin

  process_and_or : process(a,b,d,e) is

  begin

  end process process_and_or;

  process_and_or : postponed process(a,b,d,e) is

  begin

  end postponed process process_and_or;

  process_and_or : postponed process is
  begin
  end postponed process process_and_or;

  process_and_or : postponed process
  begin
  end postponed process process_and_or;

  process_and_or : process
  begin
  end process process_and_or;

  process
  begin
  end process;

  process is
  begin
  end process;

end architecture RTL;
