
architecture RTL of FIFO is

  function func_1 (a : integer) return integer is
    constant c : integer;
    variable v : integer;
    file f     : something;
  begin
  end function func1;

  function func_1 (a : integer) return integer is
    constant c   : integer;
    variable v : integer;
    file f         : something;
  begin
  end function func1;

  procedure proc_1 is
    constant c   : integer;
    variable v : integer;
    file f         : something;
  begin
  end procedure proc_1;

begin

end architecture RTL;

