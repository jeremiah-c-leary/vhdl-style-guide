
architecture RTL of FIFO is

  attribute ram_init_file : string;
  attribute ram_init_file of ram_block :
    signal is "contents.mif";


   ATTRIBUTE ram_init_file : string;

attribute      ram_init_file of ram_block :
      signal is "contents.mif";

begin

end architecture RTL;
