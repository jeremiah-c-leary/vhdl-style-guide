
architecture RTL of FIFO is

begin


  process 
  begin
  end process;

  -- Violations below

  process 
  BEGIN
  end process;

end architecture RTL;
