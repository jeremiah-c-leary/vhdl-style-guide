
context C1, C1A, C1B;

context C2, C2A, C2B;

context CON3, CON3A;
