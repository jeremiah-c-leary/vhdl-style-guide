
-- Some comment
entity FIFO is

end entity;

library ieee;

entity FIFO is

end entity;


library ieee;

-- First Comment
-- Second Comment
-- Third Comment
entity fifo is end entity;

library ieee;

-- First Comment
-- Second Comment
-- Third Comment
entity fifo is end entity;
