
entity FIFO is
BEGIN
end entity;

entity FIFO is
BEGIN
end entity;

