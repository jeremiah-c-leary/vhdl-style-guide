
architecture RTL of FIFO is

  constant c_width : integer := 16;

  CONSTANT c_depth : integer := 512;

  Constant c_word : integer := 1024;

begin

end architecture RTL;
