

architecture RTL of FIFO is

begin


end architecture RTL;
