
entity FIFO is

end entity;

entity FIFO is

end entity;

entity FIFO is

end entity;

