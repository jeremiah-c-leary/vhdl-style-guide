
library ieee;

library ieee;
