
architecture rtl of fifo is

  constant con_1 : natural := 20e10;
  constant con_2 : natural := 20.56e10;
  constant con_3 : natural := 20e-10;
  constant con_4 : natural := 20.56e-10;

  constant con_5 : natural := 20e10;
  constant con_6 : natural := 20.56e10;
  constant con_7 : natural := 20e-10;
  constant con_8 : natural := 20.56e-10;

begin

end architecture rtl;
