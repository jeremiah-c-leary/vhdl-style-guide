
architecture RTL of FIFO is

  type Voltage_Level is range 0 to 5;

  type Int_64K is range -65536 to 65535;

  type WORD is range 31 downto 0;

begin

end architecture RTL;
