
architecture rtl of fifo is

  type t_record is record
    a : std_logic;
    b : std_logic;
  end record t_record;

  type t_record is record
    a : std_logic;
    b : std_logic;
  end record t_record
  ;

  type t_record is record a : std_logic; b : std_logic; end record
  ;

  type my_array1 is array (natural range 0 to 3) of std_logic ;   -- white space before semicolon here

begin

end architecture rtl;
