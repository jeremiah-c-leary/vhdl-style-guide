
entity FIFO is

end entity FIFO;

package my_pkg is

end package my_pkg;

-- Violation below

entity FIFO is

end entity FIFO;
package my_pkg is

end package my_pkg;

