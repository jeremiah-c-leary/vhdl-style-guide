
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  PROCEDURE PROC1 IS BEGIN end PROCEDURE PROC1;

  function func1 return integer is begin End function func1;

begin

end architecture RTL;
