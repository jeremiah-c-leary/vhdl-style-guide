package test is

  type flag_pt is protected
  end protected;

  type flag_pt is protected
  end PROTECTED;

end package test;

architecture rtl of test is

  type flag_pt is protected
  end protected;

  type flag_pt is protected
  end PROTECTED;

begin

end architecture rtl;
