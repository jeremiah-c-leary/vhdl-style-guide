
architecture RTL of FIFO is

begin


  process 
  begin
  end process;

  -- Violations below

  PROCESS 
  begin
  end process;

end architecture RTL;
