

package PACK_NAME is

end package PACK_NAME;

package body PACK_NAME is

end PACK_NAME;

