
architecture RTL of FIFO is

  ATTRIBUTE max_delay : time;

  ATTRIBUTE MAX_DELAY : TIME;

begin

end architecture RTL;
