
LIBRARY ieee;

LIBRARY ieee;
