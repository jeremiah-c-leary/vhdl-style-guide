
architecture rtl of fifo is

  procedure proc is
  begin
  end;

  procedure proc is
  begin
  end;

  function func return integer is
  begin
  end func;

  function func return integer is
  begin
  end;

  procedure proc;

  function func return integer is
  begin
  end;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end;

  procedure proc is

    function func return integer is
    begin
    end func;

  begin
  end;

begin

end architecture rtl;
