
architecture RTL of ENT is
BEGIN
end RTL;

architecture RTL of ENT is
BEGIN
end rtl;

architecture RTL of ENT is
BEGIN
end Rtl;

architecture RTL of ENT is
BEGIN
end;

architecture RTL of ENT is
BEGIN
end architecture;

