
--This should pass
context con1 IS

end context con1;

--These should fail
context con1 IS
end context con1;

context co1 IS

end context con1;
