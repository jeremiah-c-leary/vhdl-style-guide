
architecture RTL of FIFO is

  attribute max_delay : time;

  ATTRIBUTE MAX_DELAY : time;

begin

end architecture RTL;
