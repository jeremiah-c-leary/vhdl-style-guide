
entity FIFO is

end entity;


entity FIFO --Comment
--Comment
--Comment
 is

end entity;
