
architecture RTL of FIFO is

  type memory is array (natural range<>) of std_logic_vector(3 downto 0);

  type memory is array (natural range<>, natural range <>) of std_logic_vector(3 downto 0);

begin

end architecture RTL;
