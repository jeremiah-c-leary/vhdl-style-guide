architecture rtl of fifo is

  signal rd_en : std_logic;
  signal wr_en : std_logic;

begin

end architecture rtl;

architecture rtl of fifo is

  signal rd_en:std_logic;
  signal wr_en:std_logic;

begin

end  architecture rtl;

architecture rtl of fifo is

  signal rd_en    :        std_logic;
  signal wr_en    :        std_logic;

begin

end  architecture rtl;
