
architecture rtl of fifo is

  -- Type attributes
  signal a : something'Ascending;
  signal a : something'Base;
  signal a : something'High;
  signal a : something'Image(x);
  signal a : something'Left;
  signal a : something'LeftOf(x);
  signal a : something'Low;
  signal a : something'Pos(x);
  signal a : something'Pred(x);
  signal a : something'Right;
  signal a : something'RightOf(x);
  signal a : something'Succ(x);
  signal a : something'Val(x);
  signal a : something'Value(x);

  -- Array attributes
  signal a : something'Ascending(n);
  signal a : something'High(n);
  signal a : something'Left(n);
  signal a : something'Length(n);
  signal a : something'Low(n);
  signal a : something'Range(n);
  signal a : something'Reverse_Range(n);
  signal a : something'Right(n);

  -- Signal attributes
  signal a : something'Active;
  signal a : something'Delayed(t);
  signal a : something'Driving;
  signal a : something'Driving_value;
  signal a : something'Event;
  signal a : something'Last_Event;
  signal a : something'Last_Active;
  signal a : something'Last_Value;
  signal a : something'Quiet(t);
  signal a : something'Stable(t);
  signal a : something'Transaction;

  -- Other attributes
  signal a : something'Instance_Name;
  signal a : something'Path_Name;
  signal a : something'Simple_name;

begin

end architecture rtl;
