
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--+-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--!-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--!---------------------------------[ abcdef ]==================================
-- Comment
--------------------------------------------------------------------------------

--!-[ abcdef ]==================================================================
-- Comment
--------------------------------------------------------------------------------

--!------------------------------------------------------------------[ abcdef ]=
-- Comment
--------------------------------------------------------------------------------

-- comment
-- comment
