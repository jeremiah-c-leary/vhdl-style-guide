
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate
    WHEN choice =>

  end generate;

  GEN_LABEL : case expression generate
    WHEN choice =>

  end generate;

end architecture;
