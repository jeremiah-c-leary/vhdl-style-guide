
architecture rtl of fifo is

  -- synthesis translate_off
  component my_block is
  end component;


  -- synthesis translate_off

  component my_block is
  end component;

begin

end architecture;
