
architecture RTL of FIFO is

begin


  process 
  begin
  end process;

  -- Violations below

  process 
  begin
  end PROCESS;

end architecture RTL;
