
architecture rtl of fifo is

begin

  PROC_LABEL : process begin end process;

  PROC_LABEL: process begin end process;

  -- Comment
PROC_LABEL : process begin end process;

  -- Comment



PROC_LABEL : process begin end process;

end;
