

library ieee;

library ieee, lib2, lib3;


