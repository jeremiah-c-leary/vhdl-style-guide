
-- Some comment
entity FIFO is

end entity;

library ieee;

entity FIFO is

end entity;

