
package body FIFO_PKG is

end package body fifo_pkg;

package body FIFO_PKG is

end package body fifo_pkg;

