
architecture rtl of fifo is

begin

  process begin

    loop end loop;

    LOOP end LOOP;

  end process;

end;
