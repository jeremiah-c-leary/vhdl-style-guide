
architecture RTL of FIFO is

begin


  process 
  begin
  end process;

  -- Violations below

  process 
  begin
  END process;

end architecture RTL;
