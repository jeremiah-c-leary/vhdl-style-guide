
package fifo_pkg is

  signal sig1 : std_logic;

end package;

package fifo_pkg is
  signal sig1 : std_logic;

end package;

