
package fifo_pkg is

end package;

package FIFO_PKG is

end package;
