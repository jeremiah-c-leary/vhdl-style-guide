

use ieee.std_logic_1164.all;

use My_Lib, OtherLib.my_math_stuff.multiply;

use YetAnotherLib.std_logic;

