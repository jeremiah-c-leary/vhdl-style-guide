
entity fifo is

end entity;

entity fifo is

end entity;

entity fifo is

end entity;

entity my_fifo is

end entity;

entity my_fifo is

end entity;

entity myfifo is

end entity;

entity myfifo is

end entity;

