
architecture rtl of fifo is

  type integer_file is file of integer;

  type integer_file is FILE of integer;

  type integer_file is File of integer;

begin

end;
