
architecture RTL of FIFO is

  signal sig1, sig2 : std_logic;
  signal sig2, sig3 : std_logic;



  signal signal1a, signal1b : std_logic;
  signal sig2a, sig2b : std_logic;


begin

end architecture RTL;
