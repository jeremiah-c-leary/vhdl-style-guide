
architecture ARCH of ENTITY is

begin

  process (one, two, three) is
  begin

  end process;

  process (one, two,
           three) is
  begin

  end  process;

  process (one, two,
           three
          ) is
  begin

  end  process;

  process (one,
           two,
           three) is
  begin

  end  process;

  process (one,
           two,
           three
          ) is
  begin

  end  process;
  process (one,
           two, three) is
  begin

  end  process;

  process (one,
           two, three
          ) is
  begin

  end  process;

  process (one, two,
           three,
           four) is
  begin

  end  process;

  process (one) is
  begin

  end  process;

  process (one
          ) is
  begin

  end  process;

  process (
           one
          ) is
  begin

  end  process;

  process (one,
           two, three,
           four,
           five, six, seven,
           eight) is
  begin

  end  process;


end architecture ARCH;

