
architecture RTL of ENT is
begin
end;

ARCHITECTURE RTL of ENT is
begin
END;

ArChItEcTuRe RTL of ENT is
begin
End;
