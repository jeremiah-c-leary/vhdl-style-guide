 
	library ieee;

library	ieee;

library 	 ieee;    
   
library 	ieee;	

library	 ieee;


-- Comment	with tab

-- Comment 	with tab

-- Comment	 with tab

-- Comment 	 with tab

-- Comment with tab	

-- Comment with tab 	

-- Comment with tab	 
