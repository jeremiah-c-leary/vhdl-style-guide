architecture rtl of fifo is

  signal sig8 : blah std_logic_vector(open);
  signal sig8 : blah std_logic_vector(37 downto 0);
  signal sig8 : blah std_logic_vector(37 downto 0, 56 downto 32);
  signal sig8 : blah std_logic_vector(37 downto 0, 56 downto 32)(5 downto 0);

  signal sig8 : std_logic_vector(open);
  signal sig8 : std_logic_vector(37 downto 0);
  signal sig8 : std_logic_vector(37 downto 0, 56 downto 32);
  signal sig8 : std_logic_vector(37 downto 0, 56 downto 32)(5 downto 0);

begin

end architecture rtl;
