--
-- This should pass
--| This should pass
----------This should pass
--==================

-- This should fail
--| This should fail
----------This should pass
--
--==================


-- ¨

-- pragmas should be ignored
--vhdl_comp_off
--vhdl_comp_on

-- (2 * 4)

--! ignore Doxygen comments
--! Space required after ! for doxygen comments

--+--block comment Header
--|
--(
--*
--+--block comment footer
