
architecture rtl of fifo is

begin

  GEN_LABEL : case expression GENERATE

  end generate;

  GEN_LABEL : case expression GENERATE

  end GENERATE;

end architecture;
