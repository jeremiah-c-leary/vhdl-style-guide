

-- Comment

-- FIXME: This should trigger

-- TODO: This should trigger
