
architecture rtl of fifo is

begin

  process begin

    report    "hello";

    report "hello";

  end process;

end architecture rtl;
