

architecture ARCH of ENTITY is

  signal my_sig : t_b_array(3 downto 0)
      (
        y(7 downto 0),
        z(2 downto 0)
            (
              a(31 downto 0)
            )
      );

  signal my_sig : t_b_array(3 downto 0)
    (
      y(7 downto 0),
      z(2 downto 0)
        (
          a(31 downto 0)
        )
    );

  signal my_sig : t_b_array(3 downto 0)
 (y(7 downto 0),z(2 downto 0)
 (a(31 downto 0)));

  signal my_sig : t_b_array(3 downto 0)
 (
      y(7 downto 0),
      z(2 downto 0)
 (
          a(31 downto 0)
        )
    );

begin

end architecture ARCH;

