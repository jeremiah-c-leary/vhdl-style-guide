
package body test is

  type flag_pt is protected body
  end protected BODY;

  type flag_pt is protected body
  end protected BODY;

end package body test;

architecture rtl of test is

  type flag_pt is protected body
  end protected BODY;

  type flag_pt is protected body
  end protected BODY;

begin

end architecture rtl;
