
architecture rtl of fifo is

begin

  test1 <= REJECT 2 ns inertial 0 after 10 ns;

  test1 <= REJECT 2 ns inertial 0 after 10 ns;

end architecture;
