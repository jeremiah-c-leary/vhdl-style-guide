
architecture rtl of fifo is

  alias designator is name;

  alias DESIGNATOR is name;

begin

end architecture rtl;
