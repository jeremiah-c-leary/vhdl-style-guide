
entity FIFO is
  generic (
    G_WIDTH : integer := 256;
    G_DEPTH : integer := 32
  );
end entity FIFO;

entity FIFO is
  port (
    I_INPUT : in integer;
    O_OUTPUT : out integer
  );
end entity FIFO;


entity FIFO is
  generic (
    G_WIDTH : integer := 256;
    G_DEPTH : integer := 32
  );
end entity FIFO;

entity FIFO is
  port (
    I_INPUT : in integer;
    O_OUTPUT : out integer
  );
end entity FIFO;

