
architecture RTL of FIFO is

  procedure proc1 is
    constant   c : integer;
    variable  v  : integer;
    file     f   : something;
  begin
  end procedure proc1;

  procedure proc1 is
    constant   c : integer;
    variable  v  : integer;
    file     f   : something;
  begin
  end procedure proc1;

  function func1 return integer is
    constant   c    : integer;
    variable  v       : integer;
    file     f     : something;
  begin
  end function func1;

begin

end architecture RTL;
