library ieee;
