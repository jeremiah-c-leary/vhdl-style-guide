
context c1;

CONTEXT c2;

Context c2;
