
architecture RTL of ENTITY1 is

  subtype range_st is range 0 to 9;
  subtype width_st is range 16 to 128;

  subtype range_subt is range 0 to 9;
  subtype width_subt is range 16 to 128;

  subtype rangest is range 0 to 9;
  subtype widthst is range 16 to 128;

begin

end architecture RTL;

