architecture rtl of fifo is

  alias ident is << constant dut.test : std_logic >>;
  alias ident is << constant   dut.test : std_logic >>;
  alias ident is << constant     dut.test : std_logic >>;

  alias ident is << signal dut.test : std_logic >>;
  alias ident is << signal          dut.test : std_logic >>;
  alias ident is << signal     dut.test : std_logic >>;

  alias ident is << variable dut.test : std_logic >>;
  alias ident is << variable dut.test : std_logic >>;
  alias ident is << variable dut.test : std_logic >>;

begin

end architecture rtl;
