
entity FIFO is

end entity;

entity FIFO is

end entity;

entity FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MY_FIFO is

end entity;

entity MYFIFO is

end entity;

entity MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity E_MYFIFO is

end entity;

entity MYFIFP is

end entity;

entity MYFIFO is

end entity;

entity E_MYFIFO_A is

end entity;

entity E_MYFIFO_A is

end entity;

entity MYFIFO_A is

end entity;

entity MYFIFO_A is

end entity;

-- Test Pascal_Snake_Case

entity MYFIFO_GREENRED_BLUE is end entity;

entity E_MY_FIFO_GREEN is end entity;

entity MY_FIFO_GREEN_A is end entity;

entity E_MYFIFO_GREENRED_BLUE_A is end entity;
