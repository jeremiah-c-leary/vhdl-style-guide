
architecture rtl of fifo is

  -- synthesis translate_on
  component my_block is
  end component;


  -- synthesis translate_on
  component my_block is
  end component;

begin

end architecture;
