

use ieee.std_logic_1164.all;

use MY_LIB, OTHERLIB.my_math_stuff.multiply;

use YetAnotherLib.std_logic;

