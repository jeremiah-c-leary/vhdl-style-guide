
ENTITY FIFO is

end entity;

ENTITY FIFO is

end entity;

ENTITY FIFO is

end entity;

