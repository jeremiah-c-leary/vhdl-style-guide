
component fifo is

end component fifo;

-- Variations

component fifo is

end component;

component fifo

end component fifo;

component fifo

end component;

