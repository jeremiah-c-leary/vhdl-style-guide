
entity FIFO is

end entity;

entity FIFO is

END entity;

entity FIFO is

End entity;

