
library ieee;

library ieee;
-- Some comment
library ieee;

library ieee;

library ieee;
