
package pkg is

  procedure MY_PROC is new my_generic_proc
    generic map (
      test => 2
    );

  function MY_FUNC is new my_generic_func
    generic map (
      test => 2
    );

  procedure MY_PROC is new my_generic_proc
    generic map (
      test => 2
    );

  function MY_FUNC is new my_generic_func
    generic map (
      test => 2
    );

  procedure MY_PROC is new my_generic_proc
    generic map (
      test => 2
    );

  function MY_FUNC is new my_generic_func
    generic map (
      test => 2
    );

end package;
