
context c1 is

end context c1;

context c1 is

end context;

context c1 is

end;
