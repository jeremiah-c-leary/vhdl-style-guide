
architecture rtl of fifo is

begin

  GEN_LABEL : for x in range (3 downto 0) generate

  end generate;

  GEN_LABEL : for x in range (3 downto 0) generate

  end generate;

end architecture;
