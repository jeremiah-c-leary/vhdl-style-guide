
package test is

  type flag_pt is protected
  end PROTECTED;

  type flag_pt is protected
  end PROTECTED;

end package test;

architecture rtl of test is

  type flag_pt is protected
  end PROTECTED;

  type flag_pt is protected
  end PROTECTED;

begin

end architecture rtl;
