
architecture RTL of ENT is
begin
END;

ARCHITECTURE RTL of ENT is
begin
END;

ArChItEcTuRe RTL of ENT is
begin
END;
