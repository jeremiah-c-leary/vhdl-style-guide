
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  PROCEDURE PROC1 IS BEGIN end PROCEDURE PROC1;

begin

end architecture RTL;
