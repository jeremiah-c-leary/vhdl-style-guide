
library ieee;
 context c1, c1a, c1b;

library ieee;
 context con1;
 context con2;
 context con3;
