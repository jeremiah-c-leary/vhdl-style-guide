entity FIFO is
generic ( a : integer );
end entity FIFO;

entity FIFO is
generic (
    a : integer
);
end entity FIFO;

entity FIFO is
generic
( a : integer
)
;
end entity FIFO;
