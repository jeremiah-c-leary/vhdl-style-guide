
architecture RTL of FIFO is

  signal sig1 : std_logic;
  signal sig2 : std_logic_vector(3 DOWNTO 0);

  -- Violations below

  signal sig1 : std_logic;
  signal sig2 : std_logic_vector(3 downto 0);


begin

end architecture RTL;
