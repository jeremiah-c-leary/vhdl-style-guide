
architecture RTL of FIFO is



end architecture RTL;
