
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block is begin end block block_label;

  BLOCK_LABEL : BLOCK IS BEGIN END BLOCK BLOCK_LABEL;

end architecture RTL;
