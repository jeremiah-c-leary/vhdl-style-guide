/**

This should pass

*/

/**

This should also pass

**/
