
package fifo_pkg is

  signal wr_en        : std_logic;
  signal rd_en        : std_logic;
  constant c_constant : integer;
  alias alias1        : subtype_indicator is name;
  alias alias1        is name;

  signal wr_en        : std_logic;
  signal rd_en        : std_logic;
  constant c_constant : integer;
  alias alias1        : subtype_indicator is name;
  alias alias1        is name;

end package;
