
entity FIFO is

end;

entity FIFO is

end;

entity FIFO is

end FIFO;

entity FIFO is

end ;

entity FIFO is

end
;

entity FIFO is

end--Comment
;
