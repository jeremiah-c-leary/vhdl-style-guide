
architecture RTl of FIFO is

  component fifo is

  end component FIFO;

  -- Failures below

  component fifo is

  end component FIFO;

  component fifo is

  end component FIFO;

begin

end architecture RTL;
