entity ENTITY1 is
  port (
    I_PORT1 : in  std_logic;
    I_PORT2 : in  std_logic;

    O_PORT3 : out std_logic;
    O_PORT4 : out std_logic
  );
end entity;
