
architecture RTL OF ENT is
begin
end RTL;

architecture RTL of ent is
begin
end rtl;

architecture RTL Of Ent is
begin
end Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;

