
architecture rtl of fifo is

  alias designator is name;

  alias designator IS name;

begin

end architecture rtl;
