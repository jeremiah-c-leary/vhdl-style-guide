
architecture ARCH of ENTITY is

begin

  -- correct block format
  BLK : block is
    signal private : std_logic;
  begin
  end block BLK;

end architecture ARCH;

