
--Ignored comment

architecture RTL of FIFO is

  signal sig1 : std_logic; -- comment
  signal sig1 : std_logic; -- comment

begin

end architecture RTL;
