
package MY_PKG is new my_generic_pkg
  generic map (
    g_my_generic => 2
  );

package MY_PKG is new my_generic_pkg
  generic map (
    g_my_generic => 2
  );
