
architecture RTL of ENTITY1 is

begin

  -- Do not flag anything
  TEST : process is
  begin

  end process TEST;

end architecture RTL;
