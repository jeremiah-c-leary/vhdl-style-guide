
architecture RTL of FIFO is

  subtype STATE_MACHINE is subtype_indication;

  -- Violations below

  subtype STATE_MACHINE is subtype_indication;

begin

end architecture RTL;
