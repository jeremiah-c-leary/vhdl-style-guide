
architecture RTL of FIFO is

begin


  PROC_LABEL : process is
  begin
  end process proc_label;

  -- Violations below

  PROC_LABEL : process is
  begin
  end process proc_label;

end architecture RTL;
