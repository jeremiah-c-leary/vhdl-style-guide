
architecture RTL of FIFO is

begin

  process

  begin

    if a = '1' then
      b <= '0';
    elsif c = '1' then
      b <= '1';
    else
      if x = '1' then
        z <= '0';
      elsif x = '0' then
        z <= '1';
      else
        z <= 'Z';
      end if;
    end if;

    if a = '0' then

      case blah is

      end case;

    end if;

    -- Violations below
    if a = '1' then
      b <= '0';
    elsif c = '1' then
      b <= '1';
    else
      if x = '1' then
        z <= '0';
      elsif x = '0' then
        z <= '1';
      else
        z <= 'Z';

      end if;



    end if;

    if a = '0' then

      case blah is

      end case;




    end if;

    -- loop statements

    if a = '1' then

    elsif c = '1' then

        loop
        end loop;

    end if;

  end process;

end architecture RTL;
