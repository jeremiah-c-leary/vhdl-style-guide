
architecture RTL of FIFO is

  signal s_sig1 : std_logic;
  signal s_sig2 : std_logic;

  -- Violations below

  signal sig1 : std_logic;
  signal sig2 : std_logic;


begin

end architecture RTL;
