
architecture RTL of ENT is
begin
end RTL;

architecture RTL of ENT is
begin
end rtl;

architecture RTL of ENT is
begin
end Rtl;

architecture RTL of ENT is
begin
end;

architecture RTL of ENT is
begin
end architecture;

