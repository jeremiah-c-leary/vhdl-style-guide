
entity FIFO is

end entity FIFO;


entity --Comment
--Comment
--Comment
FIFO is

end entity FIFO
 ;

