
architecture RTL of FIFO is

  constant c_width : integer := 16;

  constant c_depth : INTEGER := 512;

  constant c_word : Integer := 1024;

begin

end architecture RTL;
