
architecture RTL of FIFO is

begin


  process
  begin
  end PROCESS;

  -- Violations below

  process
  begin
  end PROCESS;

end architecture RTL;
