
architecture ARCH of ENTITY1 is

begin

  assert boolean
    report "Something"
    severity FAILURE;

   assert boolean
  report "Something"
    severity FAILURE;


  assert boolean
   report "Something"
  severity FAILURE;

  assert boolean
  report "Something"
 severity FAILURE;

end architecture ARCH;
