
entity FIFO is

end entity FIFO;

entity FIFO is

end entity FIFO;

entity FIFO is

end entity FIFO;

