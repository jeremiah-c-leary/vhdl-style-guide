
--This should pass
CONTEXT c1 is

end context c1;

--These should fail
CONTEXT c1 is
end context c1;

CONTEXT c1 is

end context c1;
