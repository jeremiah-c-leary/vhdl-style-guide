
port ( );

port (

);

port
(
)
;
