
architecture RTL of FIFO is

begin

  IF_LABEL : if a = '1' generate

  elsif b = '1' generate

  ELSE generate

  end generate;

  -- Violations below

  IF_LABEL : if a = '1' generate

  elsif b = '1' generate

  ELSE generate

  end generate;

end;
