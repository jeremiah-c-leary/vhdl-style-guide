

architecture RTL of ENT is

begin

  -- vsg_disable_next_line process_016
  process (A) is
  begin
    -- vsg_disable_next_line process_018
  end process;

  process (A) is
  begin
  end process;

  -- vsg_disable_next_line process_016
  -- vsg_disable_next_line process_002
  process(A)is
  begin

  -- vsg_disable_next_line process_018
  end process;

  process (A) is
  begin
  end process;

  -- vsg_disable_next_line architecture_024
end architecture;
