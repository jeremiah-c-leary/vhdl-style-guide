
package fifo_pkg is

end package FIFO_PKG;

package fifo_pkg is

end package FIFO_PKG;

