
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  COMPONENT fifo is

  end component fifo;

  Component fifo is

  end component fifo;

begin

end architecture RTL;
