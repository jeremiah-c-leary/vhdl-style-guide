
--This should pass
context con1 is

end CONTEXT con1;

--These should fail
context con1 is
end CONTEXT con1;

context co1 is

end CONTEXT con1;
