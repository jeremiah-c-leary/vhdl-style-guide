
architecture RTL of FIFO is

  procedure proc1 is
  begin
  end procedure proc1;

  -- Violations follow
  procedure proc1 is
  begin
  end procedure proc1;
  procedure proc1 is
  begin
  end procedure proc1;

begin

end architecture RTL;
