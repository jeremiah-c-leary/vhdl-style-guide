
architecture RTL of FIFO is

begin

  process 
  begin
  end process;

  process (a, b)
  begin
  end process;

  process (a, b) is
  begin
  end process;

  -- Violations below

  process 
  begin
  end process;

  process (a, b)
  begin
  end process;

  process (a, b) is
  begin
  end process;

end architecture RTL;
