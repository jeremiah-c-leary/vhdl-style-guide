
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--+-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|-----------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Comment
--|--------------------------------[ abcdef ]===================================

--------------------------------------------------------------------------------
-- Comment
--|-[ abcdef ]==================================================================

--------------------------------------------------------------------------------
-- Comment
--|------------------------------------------------------------------[ abcdef ]=

architecture rtl of fifo is

  ------------------------------------------------------------------------------
  -- Comment
  --+---------------------------------------------------------------------------

begin

end architecture rtl;

-- comment
-- comment

--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment

architecture rtl of FIFO is

begin

    inst_dummy : entity lib.module
    port map (
      -- Clocks
      clk   => clk
      --
      -- Dummy comment
      --
      data_i => data_i
    );

end architecture rtl;
