
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate
    when OTHERS =>

  end generate;

  GEN_LABEL : case expression generate
    when OTHERS =>

  end generate;

end architecture;
