
architecture RTL of FIFO is

  constant C_WIDTH : integer := 16;

  constant C_DEPTH : integer := 512;

  constant C_WORD : integer := 1024;

begin

end architecture RTL;
