entity FIFO is
port ( a : integer );
end entity FIFO;

entity FIFO is
port (
    a : integer
);
end entity FIFO;

entity FIFO is
port
( a : integer
)
;
end entity FIFO;
