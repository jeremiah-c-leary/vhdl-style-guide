
use My_Math_Stuff.MY_STRING_STUFF.my_math_stuff;

use My_Math_Stuff.MY_MATH_STUFF.my_math_stuff;

use My_Logic_Stuff.MY_LOGIC_STUFF.MY_MATH_STUFF;

