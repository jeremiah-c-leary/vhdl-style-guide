
architecture rtl of fifo is

begin

  x <= a AND b OR c NAND d NOR e XOR f XNOR g;

  x <= a AND b OR c NAND d NOR e XOR f XNOR g;

end architecture;
