

library ieee;

library ieee, std, abc;

library ieee; library std; library abc;

library ieee;
  use ieee.std_logic_1164;

library ieee; use ieee.std_logic_1164; library std; use std.something.all; library abc; use abc.blah.all;

library -- COmment
ieee --comment
; --comment
use --comment
ieee.std_logic_1164.all -- comment
; --coimment

library --comment
ieee --comment
, --comment
std --comment
, --comment
abc --comment
; --comment
