
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo is

  end COMPONENT fifo;

  component fifo is

  end Component fifo;

begin

end architecture RTL;
