
library ieee;
library work;
library std;
library bad_lib;
