
architecture RTL of FIFO is

  constant c_width : integer := 16;

  constant c_depth : integer := 512;

  constant c_word : integer := 1024;

  constant zeros : std_logic_vector(31 downto 0) := (others => '0');

  constant zeros : std_logic_vector(31 downto 0) := (others => '0');

begin

end architecture RTL;
