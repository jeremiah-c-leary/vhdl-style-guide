
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate

  end generate;

  GEN_LABEL : CASE expression generate

  end generate;

end architecture;
