
architecture RTL of FIFO is

  function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
  ) return integer is
  begin
    return 0;
  end function func_name;

  pure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
  ) return integer is
  begin
    return 0;
  end function func_name;

  impure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
  ) return integer is
  begin
    return 0;
  end function func_name;

  function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
) return integer is
  begin
    return 0;
  end function func_name;

  pure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
) return integer is
  begin
    return 0;
  end function func_name;

  impure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
) return integer is
  begin
    return 0;
  end function func_name;

  function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
       ) return integer is
  begin
    return 0;
  end function func_name;

  pure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
       ) return integer is
  begin
    return 0;
  end function func_name;

  impure function func_name (
    a : integer;
    constant b : integer;
    signal c : std_logic;
    variable v : std_logic;
    file f : std_logic
       ) return integer is
  begin
    return 0;
  end function func_name;

begin

end architecture RTL;
