
architecture rtl of fifo is

  ALIAS designator is name;

  ALIAS designator is name;

begin

end architecture rtl;
