
architecture rtl of fifo is

begin

  GEN_LABEL : case expression generate

    when 1       =>
    when n_order =>
    when others  =>

  end generate;

  GEN_LABEL : CASE expression generate

    when 1       =>
    when n_order =>
    when others  =>

  end generate;

end architecture;
