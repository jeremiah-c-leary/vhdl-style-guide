
package fifo_pkg is

end package;

library ieee;

package  fifo_pkg is

end package;

-- Comment
package fifo_pkg  is

end package;
