
architecture rtl of fifo is

  alias designator_a is name;

  alias designator is name;

begin

end architecture rtl;
