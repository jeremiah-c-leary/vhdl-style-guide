
architecture RTL of FIFO is

  procedure proc1 is begin end procedure proc1;

  PROCEDURE PROC1 IS BEGIN END PROCEDURE proc1;

begin

end architecture RTL;
