
--This should pass
context CON1 is

end context CON1;

--These should fail
context con1 is
end context con1;

context Co1 is

end context Con1;
