

architecture ARCH of ent1 is

begin

  process begin

  for i in 0 to 32 loop

  end loop;

  end process;

end architecture ARCH;


