
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    return std_logic_vector(3 downto 0);

    RETURN_LABEL : return std_logic_vector(3 downto 0);

  end process;

end architecture RTL;
