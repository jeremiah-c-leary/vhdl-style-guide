
architecture RTL of FIFO is

begin

  BLOCK_LABEL : block is begin
  end block;

  BLOCK_LABEL : block is begin end block;

end architecture RTL;
