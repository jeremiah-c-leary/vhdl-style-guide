
package sample IS

  -- represents an angle in degrees (°)

  subtype my_type is natural range 0 to 365;

end package sample;
