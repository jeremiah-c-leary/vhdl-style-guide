
architecture RTl of FIFO is

  component fifo is

  end component fifo;

  -- Failures below

  component fifo is

  END component fifo;

  component fifo is

  End component fifo;

begin

end architecture RTL;
