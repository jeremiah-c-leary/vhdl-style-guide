
entity FIFO is

END entity;

entity FIFO is

END entity;

entity FIFO is

END entity;

