
architecture rtl of fifo is

  alias designator IS name;

  alias designator IS name;

begin

end architecture rtl;
