
------------------------------------------------------------------------------------------------------------------------
-- Comment
------------------------------------------------------------------------------------------------------------------------

--+-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--!-----------------------------------------------------------------------------
-- Comment
--------------------------------------------------------------------------------

--+--------------------------------[ abcdef ]===================================
-- Comment
--------------------------------------------------------------------------------

--+-[ abcdef ]==================================================================
-- Comment
--------------------------------------------------------------------------------

--+------------------------------------------------------------------[ abcdef ]=
-- Comment
--------------------------------------------------------------------------------
architecture rtl of fifo is begin
  --+-------------------------------[ abcdef ]==================================
  -- Comment
  ------------------------------------------------------------------------------
end architecture rtl;
-- comment
-- comment

--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment
--!  Doxygen comment

------------------------------<-    80 chars    ->------------------------------
--| Comment
--| Comment
--------------------------------------------------------------------------------

