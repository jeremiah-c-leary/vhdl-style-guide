
library ieee;
context name1;
use ieee.std_logic.1164;

library ieee, lib2, lib3;
context name2, name3;
use ieee.std_logic.1164, ieee.std_logic_arith.all;

library ieee, lib2, lib3;
use ieee.std_logic.1164, ieee.std_logic_arith.all;
context name4, name5, name6;
