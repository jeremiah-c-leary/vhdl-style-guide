
architecture rtl of fifo is

  subtype t_my_array is t_array      (open)(t_range);
  subtype t_my_array is t_array (open)(t_range);
  subtype t_my_array is t_array(open)(t_range);

begin

end architecture rtl;
