
architecture rtl of fifo is

begin

  process begin

    REPORT_LABEL : report "hello";

    report "hello";

  end process;

end architecture rtl;
