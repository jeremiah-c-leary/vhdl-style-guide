
architecture RTL of FIFO is

  SIGNAL sig1 : std_logic;
  SIGNAL sig2 : std_logic;

  -- Violations below

  SIGNAL sig1 : std_logic;
  SIGNAL sig2 : std_logic;


begin

end architecture RTL;
