
architecture rtl of fifo is

begin

  process begin

    loop end loop;

    loop END LOOP;

  end process;

end;
