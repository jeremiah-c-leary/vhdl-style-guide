
ARCHITECTURE RTL of ENT is
begin
end;

ARCHITECTURE RTL of ENT is
begin
end;

ARCHITECTURE RTL of ENT is
begin
end;

