
package fifo_pkg is

end fifo_pkg;

package fifo_pkg is

end fifo_pkg;

package fifo_pkg is

end;
