
architecture RTL of FIFO is

begin

  a <= b;

  BLOCK_LABEL : block is
  begin
  end block;

  a <= b;
  BLOCK_LABEL : block is
  begin
  end block;

end architecture RTL;
