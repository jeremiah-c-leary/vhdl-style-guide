library ieee;

package body fifo_pkg is

end package body;

-- Comments are allowed
package body fifo_pkg is

end package body;

-- Violation below

library ieee;
package body fifo_pkg is

end package body;
