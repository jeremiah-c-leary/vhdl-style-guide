
architecture RTL of FIFO is

  constant c_width : integer := 16;
  constant x_depth : integer := 512;
  constant word : integer := 1024;

begin

end architecture RTL;
