library work;
  use work.tb_utilities.all;
  use work.tb_wait_clock_package.all;
  use work.random_pkg.all;
  use work.dsd_types.all;
  --use work.channel_types.all;

