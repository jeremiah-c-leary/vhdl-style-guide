
architecture RTL of FIFO is

begin


  PROC_LABEL : process 
  begin
  end process;

  postponed process 
  begin
  end process;

  process 
  begin
  end process;

  -- Violations below

PROC_LABEL : process 
  begin
  end process;

     postponed process 
  begin
  end process;

   process 
  begin
  end process;

end architecture RTL;
