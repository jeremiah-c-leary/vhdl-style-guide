
     -- synthesis translate_off

architecture rtl of fifo is

--vhdl_comp_off
--vhdl_comp_on
  -- Some comment
     -- xilinx something
-- synthesis translate_off

  signal write : std_logic;

begin

end architecture rtl;
