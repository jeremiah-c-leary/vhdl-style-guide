
architecture RTL of FIFO is

  constant c_period : integer   := 20;
  signal   wr_en    : std_logic := '1';
  signal   rd_en    : std_logic := '0';
  constant c_period : std_logic := '0';

begin

end architecture RTL;

