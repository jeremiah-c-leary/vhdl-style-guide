
architecture RTL of ent is
begin
end RTL;

architecture RTL of ent is
begin
end rtl;

architecture RTL of ent is
begin
end Rtl;

architecture RTL of ent is
begin
end;

architecture RTL of ent is
begin
end architecture;
