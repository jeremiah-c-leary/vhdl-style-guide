
package fifo_pkg is

end PACKAGE;

package fifo_pkg is

end PACKAGE;

