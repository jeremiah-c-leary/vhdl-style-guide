
package body fifo_pkg is

end package body FIFO_PKG;

package body fifo_pkg is

end package body FIFO_PKG;
