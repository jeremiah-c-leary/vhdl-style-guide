
architecture RTL of FIFO is

  constant c_width : INTEGER := 16;

  constant c_depth : INTEGER := 512;

  constant c_word : INTEGER := 1024;

begin

end architecture RTL;
