
architecture RTL of ENTITY_NAME is

begin

  process
  begin

    FORCE_LABEL : sig1 <= transport a and c;

    FORCE_LABEL : sig1 <= a and c;

    sig1 <= a and c;

  end process;

end architecture RTL;
