

architecture ARCH of ENTITY is

begin

  for i in 0 to 32 loop

  end loop;

end architecture ARCH;


