
architecture RTL of ENT is begin end architecture RTL;

architecture RTL
of
ENT is
begin
end;

architecture RTL
-- Some domment
of ENT is
begin
end;

architecture RTL--some comment
of ENT is
begin
end;
