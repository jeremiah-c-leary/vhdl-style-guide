
architecture RTL of ENT is begin end architecture RTL;

architecture RTL of ENT
is
begin
end;

architecture RTL of ENT
-- Some domment
is
begin
end;

architecture RTL of ENT--some comment
is
begin
end;

