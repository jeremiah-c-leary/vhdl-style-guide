
architecture RTL of ENT is
begin
end;

ARCHITECTURE RTL of ENT is
begin
end;

ArChItEcTuRe RTL of ENT is
begin
end;
