
context c1, c1a, c1b;

context C2, C2A, C2B;

context Con3, cOn3a;
