

architecture ARCH of ENTITY is

  signal sig : std_logic_vector(31 downto 0);
   signal SIg :  std_logic_vector(31 downto 0);
  Signal sig: std_logic_vector(31 downto 0);
 signal  sig : std_logic_vector(31 downto 0);
  signal  siG : std_logic_vector(31 downto 0);
  signal sig :std_logic_vector(31 downto 0);
  siGNal sig: std_logic_vector(31 downto 0) := "0";
  signal   SIg : std_logic_vector(31 downto 0);
  signAL sig :   std_logic_vector(31 downto 0);
  signal sig :std_logic_vector(31 downto 0);
     signal sIg : std_logic_vector(31 downto 0);
  signal sig :   std_logic_vector(31 downto 0) := (others => '0');

  signal sig1, sig2 : std_logic;
  signal sig1, sig2: std_logic;
  signal sig1, sig2 :std_logic;
  signal sig1, sig2:std_logic;

begin

end architecture ARCH;
