
architecture RTl of FIFO is

  component fifo is

  END component fifo;

  -- Failures below

  component fifo is

  END component fifo;

  component fifo is

  END component fifo;

begin

end architecture RTL;
