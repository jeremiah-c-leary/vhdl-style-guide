
architecture RTL of FIFO is

  type my_array is array(natural range <>)      of std_logic_vector(7 downto 0);
  type my_array is array(natural range <>) of std_logic_vector(7 downto 0);

begin

end architecture RTL;
