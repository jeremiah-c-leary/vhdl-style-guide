
entity FIFO is end entity;
