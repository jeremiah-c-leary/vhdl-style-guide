architecture rtl of fifo is

  variable sig8 : record_type_3(
    element1(7 downto 0),
    element2(4 downto 0)(7 downto 0)
    (
      elementA(7 downto 0),
      elementB(3 downto 0)
    ),
    element3(3 downto 0)(elementC(4 downto 1), elementD(1 downto 0)),
    element5(
      elementE
        (3 downto
            0)
        (6
 downto 0),
      elementF(7 downto 0)
    ),
    element6(4 downto
  0),
    element7(7 downto 0));

  variable sig9 : t_data_struct(data(7 downto 0));

  variable sig9 : t_data_struct(
    data(7 downto 0)
  );

begin

end architecture rtl;
