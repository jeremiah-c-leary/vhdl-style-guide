
architecture RTL of FIFO is

begin

  FOR_LABEL : for i in 0 to 7 generate

  END generate;

  IF_LABEL : if a = '1' generate

  END generate;

  CASE_LABEL : case data generate

  END generate;

  -- Violations below

  FOR_LABEL : for i in 0 to 7 generate

  END generate;

  IF_LABEL : if a = '1' generate

  END generate;

  CASE_LABEL : case data generate

  END generate;

end;
