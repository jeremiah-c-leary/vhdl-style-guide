
library ieee;
  USE ieee.std_logic_1164.all;

library ieee;
  USE ieee.std_logic_1164.all;
