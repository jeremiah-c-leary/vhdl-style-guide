 
library ieee;

library ieee;  --comment

-- Violations below

library ieee;    
   
library ieee;  -- comment      

library ieee;  -- comment      

library ieee;	

library ieee; 	

library ieee;	 

-- Comment	

-- Comment	 

-- Comment	 

