
architecture RTL of FIFO is

  FILE defaultImage : load_file_type open read_mode is load_file_name;

  FILE defaultImage : load_file_type open read_mode is load_file_name;

  FILE defaultImage : load_file_type open read_mode is load_file_name;

begin

end;
