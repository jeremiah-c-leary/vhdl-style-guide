
architecture rtl of fifo is

begin

  gen_label : for x IN range (3 downto 0) generate

  end generate;

  gen_label : for x IN range (3 downto 0) generate

  end generate;

end architecture;
