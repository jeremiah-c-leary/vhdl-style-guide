
architecture RTL of FIFO is

  constant width_c : integer := 16;
  constant depth_x : integer := 512;
  constant word : integer := 1024;

begin

end architecture RTL;
