

library lib1;
-- Comment 1
  use lib1.all;

library lib2;
  -- Comment 2
  use lib2.all;

