
architecture rtl of fifo is

  file defaultimage : load_file_type open read_mode IS load_file_name;

  file defaultimage : load_file_type open read_mode IS load_file_name;

  file defaultimage : load_file_type open read_mode IS load_file_name;

begin

end;
