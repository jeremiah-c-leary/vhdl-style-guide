
architecture RTL of FIFO is

  subtype state_machine is subtype_indication;

  -- Violations below

  SUBTYPE state_machine is subtype_indication;

begin

end architecture RTL;
